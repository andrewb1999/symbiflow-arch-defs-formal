module top(
  input clk,
  input [7:0] sw,
  output [7:0] led
  );
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A1;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A2;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A3;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A4;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_AO5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_AO6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_AQ;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_AX;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A_CY;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A_XOR;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B1;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B2;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B3;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B4;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_BMUX;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_BO5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_BO6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_BQ;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_BX;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B_CY;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B_XOR;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C1;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C2;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C3;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C4;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_CLK;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_CMUX;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_CO5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_CO6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_COUT;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_CQ;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_CX;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C_CY;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C_XOR;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D1;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D2;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D3;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D4;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_DMUX;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_DO5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_DO6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_DQ;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_DX;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D_CY;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D_XOR;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A1;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A2;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A3;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A4;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_AO5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_AO6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A_CY;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A_XOR;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B1;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B2;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B3;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B4;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_BO5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_BO6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B_CY;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B_XOR;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C1;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C2;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C3;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C4;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_CO5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_CO6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C_CY;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C_XOR;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D1;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D2;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D3;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D4;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_DO5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_DO6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D_CY;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D_XOR;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A1;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A2;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A3;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A4;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_AMUX;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_AO5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_AO6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_AQ;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_AX;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A_CY;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A_XOR;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B1;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B2;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B3;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B4;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_BMUX;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_BO5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_BO6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_BQ;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_BX;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B_CY;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B_XOR;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C1;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C2;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C3;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C4;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_CIN;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_CLK;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_CMUX;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_CO5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_CO6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_COUT;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_CQ;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_CX;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C_CY;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C_XOR;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D1;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D2;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D3;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D4;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_DMUX;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_DO5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_DO6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_DQ;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_DX;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D_CY;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D_XOR;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A1;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A2;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A3;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A4;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_AO5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_AO6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A_CY;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A_XOR;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B1;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B2;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B3;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B4;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_BO5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_BO6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B_CY;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B_XOR;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C1;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C2;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C3;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C4;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_CO5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_CO6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C_CY;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C_XOR;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D1;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D2;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D3;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D4;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_DO5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_DO6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D_CY;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D_XOR;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_A;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_A1;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_A2;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_A3;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_A4;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_A5;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_A6;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_AMUX;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_AO5;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_AO6;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_AQ;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_AX;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_A_CY;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_A_XOR;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_B;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_B1;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_B2;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_B3;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_B4;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_B5;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_B6;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_BMUX;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_BO5;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_BO6;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_BQ;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_BX;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_B_CY;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_B_XOR;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_C;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_C1;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_C2;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_C3;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_C4;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_C5;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_C6;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_CIN;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_CLK;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_CMUX;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_CO5;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_CO6;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_COUT;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_CQ;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_CX;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_C_CY;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_C_XOR;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_D;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_D1;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_D2;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_D3;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_D4;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_D5;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_D6;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_DMUX;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_DO5;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_DO6;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_DQ;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_DX;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_D_CY;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X26Y127_D_XOR;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_A;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_A1;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_A2;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_A3;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_A4;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_A5;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_A6;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_AO5;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_AO6;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_A_CY;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_A_XOR;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_B;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_B1;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_B2;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_B3;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_B4;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_B5;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_B6;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_BO5;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_BO6;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_B_CY;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_B_XOR;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_C;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_C1;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_C2;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_C3;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_C4;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_C5;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_C6;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_CO5;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_CO6;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_C_CY;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_C_XOR;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_D;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_D1;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_D2;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_D3;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_D4;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_D5;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_D6;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_DO5;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_DO6;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_D_CY;
  wire [0:0] CLBLL_R_X17Y127_SLICE_X27Y127_D_XOR;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A1;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A2;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A3;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A4;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_AMUX;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_AO5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_AO6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_AQ;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_AX;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A_CY;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A_XOR;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B1;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B2;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B3;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B4;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_BMUX;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_BO5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_BO6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_BQ;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_BX;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B_CY;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B_XOR;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C1;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C2;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C3;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C4;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_CIN;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_CLK;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_CMUX;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_CO5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_CO6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_COUT;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_CQ;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_CX;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C_CY;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C_XOR;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D1;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D2;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D3;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D4;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_DMUX;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_DO5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_DO6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_DQ;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_DX;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D_CY;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D_XOR;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A1;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A2;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A3;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A4;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_AO5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_AO6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A_CY;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A_XOR;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B1;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B2;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B3;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B4;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_BO5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_BO6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B_CY;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B_XOR;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C1;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C2;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C3;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C4;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_CO5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_CO6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C_CY;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C_XOR;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D1;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D2;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D3;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D4;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_DO5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_DO6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D_CY;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D_XOR;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A1;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A2;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A3;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A4;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_AO5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_AO6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_AQ;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_AX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A_CY;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A_XOR;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B1;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B2;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B3;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B4;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_BMUX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_BO5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_BO6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_BQ;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_BX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B_CY;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B_XOR;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C1;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C2;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C3;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C4;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_CIN;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_CLK;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_CMUX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_CO5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_CO6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_COUT;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_CQ;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_CX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C_CY;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C_XOR;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D1;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D2;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D3;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D4;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_DMUX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_DO5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_DO6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_DQ;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_DX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D_CY;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D_XOR;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A1;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A2;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A3;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A4;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_AO5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_AO6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A_CY;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A_XOR;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B1;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B2;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B3;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B4;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_BO5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_BO6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B_CY;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B_XOR;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C1;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C2;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C3;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C4;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_CO5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_CO6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C_CY;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C_XOR;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D1;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D2;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D3;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D4;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_DO5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_DO6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D_CY;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D_XOR;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A1;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A2;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A3;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A4;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_AO5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_AO6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_AQ;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_AX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A_CY;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A_XOR;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B1;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B2;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B3;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B4;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_BMUX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_BO5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_BO6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_BQ;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_BX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B_CY;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B_XOR;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C1;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C2;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C3;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C4;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_CIN;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_CLK;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_CMUX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_CO5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_CO6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_COUT;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_CQ;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_CX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C_CY;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C_XOR;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D1;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D2;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D3;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D4;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_DMUX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_DO5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_DO6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_DQ;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_DX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D_CY;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D_XOR;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A1;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A2;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A3;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A4;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_AO5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_AO6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A_CY;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A_XOR;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B1;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B2;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B3;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B4;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_BO5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_BO6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B_CY;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B_XOR;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C1;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C2;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C3;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C4;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_CO5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_CO6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C_CY;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C_XOR;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D1;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D2;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D3;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D4;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_DO5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_DO6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D_CY;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D_XOR;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A1;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A2;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A3;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A4;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_AO5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_AO6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_AQ;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_AX;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A_CY;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A_XOR;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B1;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B2;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B3;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B4;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_BMUX;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_BO5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_BO6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_BQ;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_BX;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B_CY;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B_XOR;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C1;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C2;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C3;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C4;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_CIN;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_CLK;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_CMUX;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_CO5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_CO6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_COUT;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_CQ;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_CX;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C_CY;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C_XOR;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D1;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D2;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D3;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D4;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_DMUX;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_DO5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_DO6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_DQ;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_DX;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D_CY;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D_XOR;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A1;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A2;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A3;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A4;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_AO5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_AO6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A_CY;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A_XOR;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B1;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B2;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B3;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B4;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_BO5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_BO6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B_CY;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B_XOR;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C1;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C2;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C3;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C4;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_CO5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_CO6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C_CY;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C_XOR;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D1;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D2;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D3;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D4;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_DO5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_DO6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D_CY;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D_XOR;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A1;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A2;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A3;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A4;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_AO5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_AO6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_AQ;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_AX;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A_CY;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A_XOR;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B1;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B2;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B3;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B4;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_BMUX;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_BO5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_BO6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_BQ;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_BX;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B_CY;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B_XOR;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C1;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C2;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C3;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C4;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_CIN;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_CLK;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_CMUX;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_CO5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_CO6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_COUT;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_CQ;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_CX;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C_CY;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C_XOR;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D1;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D2;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D3;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D4;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_DMUX;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_DO5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_DO6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_DQ;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_DX;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D_CY;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D_XOR;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A1;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A2;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A3;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A4;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_AO5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_AO6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A_CY;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A_XOR;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B1;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B2;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B3;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B4;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_BO5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_BO6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B_CY;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B_XOR;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C1;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C2;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C3;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C4;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_CO5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_CO6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C_CY;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C_XOR;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D1;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D2;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D3;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D4;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_DO5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_DO6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D_CY;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D_XOR;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_A;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_A1;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_A2;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_A3;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_A4;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_A5;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_A6;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_AO5;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_AO6;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_AQ;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_AX;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_A_CY;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_A_XOR;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_B;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_B1;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_B2;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_B3;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_B4;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_B5;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_B6;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_BMUX;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_BO5;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_BO6;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_BQ;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_BX;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_B_CY;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_B_XOR;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_C;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_C1;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_C2;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_C3;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_C4;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_C5;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_C6;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_CIN;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_CLK;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_CMUX;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_CO5;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_CO6;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_COUT;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_CQ;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_CX;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_C_CY;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_C_XOR;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_D;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_D1;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_D2;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_D3;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_D4;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_D5;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_D6;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_DMUX;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_DO5;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_DO6;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_DQ;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_DX;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_D_CY;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X26Y133_D_XOR;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_A;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_A1;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_A2;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_A3;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_A4;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_A5;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_A6;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_AO5;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_AO6;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_A_CY;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_A_XOR;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_B;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_B1;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_B2;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_B3;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_B4;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_B5;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_B6;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_BO5;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_BO6;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_B_CY;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_B_XOR;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_C;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_C1;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_C2;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_C3;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_C4;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_C5;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_C6;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_CO5;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_CO6;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_C_CY;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_C_XOR;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_D;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_D1;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_D2;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_D3;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_D4;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_D5;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_D6;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_DO5;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_DO6;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_D_CY;
  wire [0:0] CLBLL_R_X17Y133_SLICE_X27Y133_D_XOR;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S1;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_CE;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_I;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_I;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_O;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y2_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_TQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_TQ;
  wire [0:0] RIOB33_SING_X43Y50_IOB_X1Y50_O;
  wire [0:0] RIOB33_X43Y51_IOB_X1Y51_O;
  wire [0:0] RIOB33_X43Y51_IOB_X1Y52_O;
  wire [0:0] RIOB33_X43Y55_IOB_X1Y55_O;
  wire [0:0] RIOB33_X43Y57_IOB_X1Y58_O;
  wire [0:0] RIOB33_X43Y61_IOB_X1Y61_O;
  wire [0:0] RIOB33_X43Y75_IOB_X1Y76_I;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_D1;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_OQ;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_T1;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_TQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_D1;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_OQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_T1;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_TQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_D1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_OQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_T1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_TQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_D1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_OQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_T1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_TQ;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_D1;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_OQ;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_T1;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_TQ;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_D1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_OQ;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_T1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_TQ;
  wire [0:0] RIOI3_X43Y75_ILOGIC_X1Y76_D;
  wire [0:0] RIOI3_X43Y75_ILOGIC_X1Y76_O;
  wire [0:0] \$abc$3569$aiger3568$100 ;
  wire [0:0] \$abc$3569$aiger3568$109 ;
  wire [0:0] \$abc$3569$aiger3568$118 ;
  wire [0:0] \$abc$3569$aiger3568$55 ;
  wire [0:0] \$abc$3569$aiger3568$64 ;
  wire [0:0] \$abc$3569$aiger3568$73 ;
  wire [0:0] \$abc$3569$aiger3568$82 ;
  wire [0:0] \$abc$3569$aiger3568$91 ;
  wire [35:0] \$auto$alumacc.cc:485:replace_alu$1385.O ;
  wire [27:0] \counter ;


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1471CLBLL_R_X17Y125_SLICE_X26Y125_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y125_SLICE_X26Y125_AO6),
.Q(\counter [0]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1473CLBLL_R_X17Y125_SLICE_X26Y125_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y125_SLICE_X26Y125_BO5),
.Q(\counter [2]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1474CLBLL_R_X17Y125_SLICE_X26Y125_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y125_SLICE_X26Y125_CO5),
.Q(\counter [3]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1472CLBLL_R_X17Y125_SLICE_X26Y125_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y125_SLICE_X26Y125_DO5),
.Q(\counter [1]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y125_SLICE_X26Y125_CARRY4 (
.CI(1'b0),
.CO({\$abc$3569$aiger3568$55 , CLBLL_R_X17Y125_SLICE_X26Y125_C_CY, CLBLL_R_X17Y125_SLICE_X26Y125_B_CY, CLBLL_R_X17Y125_SLICE_X26Y125_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({\$auto$alumacc.cc:485:replace_alu$1385.O [3], \$auto$alumacc.cc:485:replace_alu$1385.O [2], \$auto$alumacc.cc:485:replace_alu$1385.O [1], CLBLL_R_X17Y125_SLICE_X26Y125_A_XOR}),
.S({CLBLL_R_X17Y125_SLICE_X26Y125_DO6, CLBLL_R_X17Y125_SLICE_X26Y125_CO6, CLBLL_R_X17Y125_SLICE_X26Y125_BO6, CLBLL_R_X17Y125_SLICE_X26Y125_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff00ff00)
  ) CLBLL_R_X17Y125_SLICE_X26Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(\$auto$alumacc.cc:485:replace_alu$1385.O [1]),
.I4(\counter [3]),
.I5(1'b1),
.O5(CLBLL_R_X17Y125_SLICE_X26Y125_DO5),
.O6(CLBLL_R_X17Y125_SLICE_X26Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaaaaaaa)
  ) CLBLL_R_X17Y125_SLICE_X26Y125_CLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1385.O [3]),
.I1(1'b1),
.I2(\counter [2]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y125_SLICE_X26Y125_CO5),
.O6(CLBLL_R_X17Y125_SLICE_X26Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0f0f0f0)
  ) CLBLL_R_X17Y125_SLICE_X26Y125_BLUT (
.I0(1'b1),
.I1(\counter [1]),
.I2(\$auto$alumacc.cc:485:replace_alu$1385.O [2]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y125_SLICE_X26Y125_BO5),
.O6(CLBLL_R_X17Y125_SLICE_X26Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00000000)
  ) CLBLL_R_X17Y125_SLICE_X26Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(\counter [0]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y125_SLICE_X26Y125_AO5),
.O6(CLBLL_R_X17Y125_SLICE_X26Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y125_SLICE_X27Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y125_SLICE_X27Y125_DO5),
.O6(CLBLL_R_X17Y125_SLICE_X27Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y125_SLICE_X27Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y125_SLICE_X27Y125_CO5),
.O6(CLBLL_R_X17Y125_SLICE_X27Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y125_SLICE_X27Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y125_SLICE_X27Y125_BO5),
.O6(CLBLL_R_X17Y125_SLICE_X27Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y125_SLICE_X27Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y125_SLICE_X27Y125_AO5),
.O6(CLBLL_R_X17Y125_SLICE_X27Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1477CLBLL_R_X17Y126_SLICE_X26Y126_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y126_SLICE_X26Y126_AO5),
.Q(\counter [6]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1478CLBLL_R_X17Y126_SLICE_X26Y126_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y126_SLICE_X26Y126_BO5),
.Q(\counter [7]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1475CLBLL_R_X17Y126_SLICE_X26Y126_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y126_SLICE_X26Y126_CO5),
.Q(\counter [4]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1476CLBLL_R_X17Y126_SLICE_X26Y126_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y126_SLICE_X26Y126_DO5),
.Q(\counter [5]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y126_SLICE_X26Y126_CARRY4 (
.CI(\$abc$3569$aiger3568$55 ),
.CO({\$abc$3569$aiger3568$64 , CLBLL_R_X17Y126_SLICE_X26Y126_C_CY, CLBLL_R_X17Y126_SLICE_X26Y126_B_CY, CLBLL_R_X17Y126_SLICE_X26Y126_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1385.O [7], \$auto$alumacc.cc:485:replace_alu$1385.O [6], \$auto$alumacc.cc:485:replace_alu$1385.O [5], \$auto$alumacc.cc:485:replace_alu$1385.O [4]}),
.S({CLBLL_R_X17Y126_SLICE_X26Y126_DO6, CLBLL_R_X17Y126_SLICE_X26Y126_CO6, CLBLL_R_X17Y126_SLICE_X26Y126_BO6, CLBLL_R_X17Y126_SLICE_X26Y126_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLL_R_X17Y126_SLICE_X26Y126_DLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1385.O [5]),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(\counter [7]),
.I5(1'b1),
.O5(CLBLL_R_X17Y126_SLICE_X26Y126_DO5),
.O6(CLBLL_R_X17Y126_SLICE_X26Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_R_X17Y126_SLICE_X26Y126_CLUT (
.I0(1'b1),
.I1(\$auto$alumacc.cc:485:replace_alu$1385.O [4]),
.I2(\counter [6]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y126_SLICE_X26Y126_CO5),
.O6(CLBLL_R_X17Y126_SLICE_X26Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y126_SLICE_X26Y126_BLUT (
.I0(1'b1),
.I1(\counter [5]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1385.O [7]),
.I5(1'b1),
.O5(CLBLL_R_X17Y126_SLICE_X26Y126_BO5),
.O6(CLBLL_R_X17Y126_SLICE_X26Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y126_SLICE_X26Y126_ALUT (
.I0(1'b1),
.I1(\counter [4]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1385.O [6]),
.I5(1'b1),
.O5(CLBLL_R_X17Y126_SLICE_X26Y126_AO5),
.O6(CLBLL_R_X17Y126_SLICE_X26Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y126_SLICE_X27Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y126_SLICE_X27Y126_DO5),
.O6(CLBLL_R_X17Y126_SLICE_X27Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y126_SLICE_X27Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y126_SLICE_X27Y126_CO5),
.O6(CLBLL_R_X17Y126_SLICE_X27Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y126_SLICE_X27Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y126_SLICE_X27Y126_BO5),
.O6(CLBLL_R_X17Y126_SLICE_X27Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y126_SLICE_X27Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y126_SLICE_X27Y126_AO5),
.O6(CLBLL_R_X17Y126_SLICE_X27Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1481CLBLL_R_X17Y127_SLICE_X26Y127_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y127_SLICE_X26Y127_AO5),
.Q(\counter [10]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1482CLBLL_R_X17Y127_SLICE_X26Y127_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y127_SLICE_X26Y127_BO5),
.Q(\counter [11]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1479CLBLL_R_X17Y127_SLICE_X26Y127_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y127_SLICE_X26Y127_CO5),
.Q(\counter [8]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1480CLBLL_R_X17Y127_SLICE_X26Y127_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y127_SLICE_X26Y127_DO5),
.Q(\counter [9]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y127_SLICE_X26Y127_CARRY4 (
.CI(\$abc$3569$aiger3568$64 ),
.CO({\$abc$3569$aiger3568$73 , CLBLL_R_X17Y127_SLICE_X26Y127_C_CY, CLBLL_R_X17Y127_SLICE_X26Y127_B_CY, CLBLL_R_X17Y127_SLICE_X26Y127_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1385.O [11], \$auto$alumacc.cc:485:replace_alu$1385.O [10], \$auto$alumacc.cc:485:replace_alu$1385.O [9], \$auto$alumacc.cc:485:replace_alu$1385.O [8]}),
.S({CLBLL_R_X17Y127_SLICE_X26Y127_DO6, CLBLL_R_X17Y127_SLICE_X26Y127_CO6, CLBLL_R_X17Y127_SLICE_X26Y127_BO6, CLBLL_R_X17Y127_SLICE_X26Y127_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLL_R_X17Y127_SLICE_X26Y127_DLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1385.O [9]),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(\counter [11]),
.I5(1'b1),
.O5(CLBLL_R_X17Y127_SLICE_X26Y127_DO5),
.O6(CLBLL_R_X17Y127_SLICE_X26Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_R_X17Y127_SLICE_X26Y127_CLUT (
.I0(1'b1),
.I1(\$auto$alumacc.cc:485:replace_alu$1385.O [8]),
.I2(\counter [10]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y127_SLICE_X26Y127_CO5),
.O6(CLBLL_R_X17Y127_SLICE_X26Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y127_SLICE_X26Y127_BLUT (
.I0(1'b1),
.I1(\counter [9]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1385.O [11]),
.I5(1'b1),
.O5(CLBLL_R_X17Y127_SLICE_X26Y127_BO5),
.O6(CLBLL_R_X17Y127_SLICE_X26Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y127_SLICE_X26Y127_ALUT (
.I0(1'b1),
.I1(\counter [8]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1385.O [10]),
.I5(1'b1),
.O5(CLBLL_R_X17Y127_SLICE_X26Y127_AO5),
.O6(CLBLL_R_X17Y127_SLICE_X26Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y127_SLICE_X27Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y127_SLICE_X27Y127_DO5),
.O6(CLBLL_R_X17Y127_SLICE_X27Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y127_SLICE_X27Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y127_SLICE_X27Y127_CO5),
.O6(CLBLL_R_X17Y127_SLICE_X27Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y127_SLICE_X27Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y127_SLICE_X27Y127_BO5),
.O6(CLBLL_R_X17Y127_SLICE_X27Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y127_SLICE_X27Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y127_SLICE_X27Y127_AO5),
.O6(CLBLL_R_X17Y127_SLICE_X27Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1485CLBLL_R_X17Y128_SLICE_X26Y128_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y128_SLICE_X26Y128_AO5),
.Q(\counter [14]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1486CLBLL_R_X17Y128_SLICE_X26Y128_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y128_SLICE_X26Y128_BO5),
.Q(\counter [15]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1483CLBLL_R_X17Y128_SLICE_X26Y128_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y128_SLICE_X26Y128_CO5),
.Q(\counter [12]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1484CLBLL_R_X17Y128_SLICE_X26Y128_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y128_SLICE_X26Y128_DO5),
.Q(\counter [13]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y128_SLICE_X26Y128_CARRY4 (
.CI(\$abc$3569$aiger3568$73 ),
.CO({\$abc$3569$aiger3568$82 , CLBLL_R_X17Y128_SLICE_X26Y128_C_CY, CLBLL_R_X17Y128_SLICE_X26Y128_B_CY, CLBLL_R_X17Y128_SLICE_X26Y128_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1385.O [15], \$auto$alumacc.cc:485:replace_alu$1385.O [14], \$auto$alumacc.cc:485:replace_alu$1385.O [13], \$auto$alumacc.cc:485:replace_alu$1385.O [12]}),
.S({CLBLL_R_X17Y128_SLICE_X26Y128_DO6, CLBLL_R_X17Y128_SLICE_X26Y128_CO6, CLBLL_R_X17Y128_SLICE_X26Y128_BO6, CLBLL_R_X17Y128_SLICE_X26Y128_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLL_R_X17Y128_SLICE_X26Y128_DLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1385.O [13]),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(\counter [15]),
.I5(1'b1),
.O5(CLBLL_R_X17Y128_SLICE_X26Y128_DO5),
.O6(CLBLL_R_X17Y128_SLICE_X26Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_R_X17Y128_SLICE_X26Y128_CLUT (
.I0(1'b1),
.I1(\$auto$alumacc.cc:485:replace_alu$1385.O [12]),
.I2(\counter [14]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y128_SLICE_X26Y128_CO5),
.O6(CLBLL_R_X17Y128_SLICE_X26Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y128_SLICE_X26Y128_BLUT (
.I0(1'b1),
.I1(\counter [13]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1385.O [15]),
.I5(1'b1),
.O5(CLBLL_R_X17Y128_SLICE_X26Y128_BO5),
.O6(CLBLL_R_X17Y128_SLICE_X26Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y128_SLICE_X26Y128_ALUT (
.I0(1'b1),
.I1(\counter [12]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1385.O [14]),
.I5(1'b1),
.O5(CLBLL_R_X17Y128_SLICE_X26Y128_AO5),
.O6(CLBLL_R_X17Y128_SLICE_X26Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y128_SLICE_X27Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y128_SLICE_X27Y128_DO5),
.O6(CLBLL_R_X17Y128_SLICE_X27Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y128_SLICE_X27Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y128_SLICE_X27Y128_CO5),
.O6(CLBLL_R_X17Y128_SLICE_X27Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y128_SLICE_X27Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y128_SLICE_X27Y128_BO5),
.O6(CLBLL_R_X17Y128_SLICE_X27Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y128_SLICE_X27Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y128_SLICE_X27Y128_AO5),
.O6(CLBLL_R_X17Y128_SLICE_X27Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1487CLBLL_R_X17Y129_SLICE_X26Y129_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y129_SLICE_X26Y129_A_XOR),
.Q(\counter [16]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1489CLBLL_R_X17Y129_SLICE_X26Y129_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y129_SLICE_X26Y129_BO5),
.Q(\counter [18]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1490CLBLL_R_X17Y129_SLICE_X26Y129_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y129_SLICE_X26Y129_CO5),
.Q(\counter [19]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1488CLBLL_R_X17Y129_SLICE_X26Y129_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y129_SLICE_X26Y129_DO5),
.Q(\counter [17]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y129_SLICE_X26Y129_CARRY4 (
.CI(\$abc$3569$aiger3568$82 ),
.CO({\$abc$3569$aiger3568$91 , CLBLL_R_X17Y129_SLICE_X26Y129_C_CY, CLBLL_R_X17Y129_SLICE_X26Y129_B_CY, CLBLL_R_X17Y129_SLICE_X26Y129_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1385.O [19], \$auto$alumacc.cc:485:replace_alu$1385.O [18], \$auto$alumacc.cc:485:replace_alu$1385.O [17], CLBLL_R_X17Y129_SLICE_X26Y129_A_XOR}),
.S({CLBLL_R_X17Y129_SLICE_X26Y129_DO6, CLBLL_R_X17Y129_SLICE_X26Y129_CO6, CLBLL_R_X17Y129_SLICE_X26Y129_BO6, CLBLL_R_X17Y129_SLICE_X26Y129_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLL_R_X17Y129_SLICE_X26Y129_DLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1385.O [17]),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(\counter [19]),
.I5(1'b1),
.O5(CLBLL_R_X17Y129_SLICE_X26Y129_DO5),
.O6(CLBLL_R_X17Y129_SLICE_X26Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_R_X17Y129_SLICE_X26Y129_CLUT (
.I0(1'b1),
.I1(\$auto$alumacc.cc:485:replace_alu$1385.O [19]),
.I2(\counter [18]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y129_SLICE_X26Y129_CO5),
.O6(CLBLL_R_X17Y129_SLICE_X26Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y129_SLICE_X26Y129_BLUT (
.I0(1'b1),
.I1(\counter [17]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1385.O [18]),
.I5(1'b1),
.O5(CLBLL_R_X17Y129_SLICE_X26Y129_BO5),
.O6(CLBLL_R_X17Y129_SLICE_X26Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLL_R_X17Y129_SLICE_X26Y129_ALUT (
.I0(1'b1),
.I1(\counter [16]),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y129_SLICE_X26Y129_AO5),
.O6(CLBLL_R_X17Y129_SLICE_X26Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y129_SLICE_X27Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y129_SLICE_X27Y129_DO5),
.O6(CLBLL_R_X17Y129_SLICE_X27Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y129_SLICE_X27Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y129_SLICE_X27Y129_CO5),
.O6(CLBLL_R_X17Y129_SLICE_X27Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y129_SLICE_X27Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y129_SLICE_X27Y129_BO5),
.O6(CLBLL_R_X17Y129_SLICE_X27Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y129_SLICE_X27Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y129_SLICE_X27Y129_AO5),
.O6(CLBLL_R_X17Y129_SLICE_X27Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1491CLBLL_R_X17Y130_SLICE_X26Y130_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y130_SLICE_X26Y130_A_XOR),
.Q(\counter [20]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1493CLBLL_R_X17Y130_SLICE_X26Y130_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y130_SLICE_X26Y130_BO5),
.Q(\counter [22]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1494CLBLL_R_X17Y130_SLICE_X26Y130_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y130_SLICE_X26Y130_CO5),
.Q(\counter [23]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1492CLBLL_R_X17Y130_SLICE_X26Y130_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y130_SLICE_X26Y130_DO5),
.Q(\counter [21]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y130_SLICE_X26Y130_CARRY4 (
.CI(\$abc$3569$aiger3568$91 ),
.CO({\$abc$3569$aiger3568$100 , CLBLL_R_X17Y130_SLICE_X26Y130_C_CY, CLBLL_R_X17Y130_SLICE_X26Y130_B_CY, CLBLL_R_X17Y130_SLICE_X26Y130_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1385.O [23], \$auto$alumacc.cc:485:replace_alu$1385.O [22], \$auto$alumacc.cc:485:replace_alu$1385.O [21], CLBLL_R_X17Y130_SLICE_X26Y130_A_XOR}),
.S({CLBLL_R_X17Y130_SLICE_X26Y130_DO6, CLBLL_R_X17Y130_SLICE_X26Y130_CO6, CLBLL_R_X17Y130_SLICE_X26Y130_BO6, CLBLL_R_X17Y130_SLICE_X26Y130_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLL_R_X17Y130_SLICE_X26Y130_DLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1385.O [21]),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(\counter [23]),
.I5(1'b1),
.O5(CLBLL_R_X17Y130_SLICE_X26Y130_DO5),
.O6(CLBLL_R_X17Y130_SLICE_X26Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_R_X17Y130_SLICE_X26Y130_CLUT (
.I0(1'b1),
.I1(\$auto$alumacc.cc:485:replace_alu$1385.O [23]),
.I2(\counter [22]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y130_SLICE_X26Y130_CO5),
.O6(CLBLL_R_X17Y130_SLICE_X26Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y130_SLICE_X26Y130_BLUT (
.I0(1'b1),
.I1(\counter [21]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1385.O [22]),
.I5(1'b1),
.O5(CLBLL_R_X17Y130_SLICE_X26Y130_BO5),
.O6(CLBLL_R_X17Y130_SLICE_X26Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLL_R_X17Y130_SLICE_X26Y130_ALUT (
.I0(1'b1),
.I1(\counter [20]),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y130_SLICE_X26Y130_AO5),
.O6(CLBLL_R_X17Y130_SLICE_X26Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y130_SLICE_X27Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y130_SLICE_X27Y130_DO5),
.O6(CLBLL_R_X17Y130_SLICE_X27Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y130_SLICE_X27Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y130_SLICE_X27Y130_CO5),
.O6(CLBLL_R_X17Y130_SLICE_X27Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y130_SLICE_X27Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y130_SLICE_X27Y130_BO5),
.O6(CLBLL_R_X17Y130_SLICE_X27Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y130_SLICE_X27Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y130_SLICE_X27Y130_AO5),
.O6(CLBLL_R_X17Y130_SLICE_X27Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1495CLBLL_R_X17Y131_SLICE_X26Y131_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y131_SLICE_X26Y131_A_XOR),
.Q(\counter [24]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1497CLBLL_R_X17Y131_SLICE_X26Y131_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y131_SLICE_X26Y131_BO5),
.Q(\counter [26]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1498CLBLL_R_X17Y131_SLICE_X26Y131_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y131_SLICE_X26Y131_CO5),
.Q(\counter [27]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1496CLBLL_R_X17Y131_SLICE_X26Y131_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y131_SLICE_X26Y131_DO5),
.Q(\counter [25]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y131_SLICE_X26Y131_CARRY4 (
.CI(\$abc$3569$aiger3568$100 ),
.CO({\$abc$3569$aiger3568$109 , CLBLL_R_X17Y131_SLICE_X26Y131_C_CY, CLBLL_R_X17Y131_SLICE_X26Y131_B_CY, CLBLL_R_X17Y131_SLICE_X26Y131_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1385.O [27], \$auto$alumacc.cc:485:replace_alu$1385.O [26], \$auto$alumacc.cc:485:replace_alu$1385.O [25], CLBLL_R_X17Y131_SLICE_X26Y131_A_XOR}),
.S({CLBLL_R_X17Y131_SLICE_X26Y131_DO6, CLBLL_R_X17Y131_SLICE_X26Y131_CO6, CLBLL_R_X17Y131_SLICE_X26Y131_BO6, CLBLL_R_X17Y131_SLICE_X26Y131_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLL_R_X17Y131_SLICE_X26Y131_DLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1385.O [25]),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(\counter [27]),
.I5(1'b1),
.O5(CLBLL_R_X17Y131_SLICE_X26Y131_DO5),
.O6(CLBLL_R_X17Y131_SLICE_X26Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_R_X17Y131_SLICE_X26Y131_CLUT (
.I0(1'b1),
.I1(\$auto$alumacc.cc:485:replace_alu$1385.O [27]),
.I2(\counter [26]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y131_SLICE_X26Y131_CO5),
.O6(CLBLL_R_X17Y131_SLICE_X26Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y131_SLICE_X26Y131_BLUT (
.I0(1'b1),
.I1(\counter [25]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1385.O [26]),
.I5(1'b1),
.O5(CLBLL_R_X17Y131_SLICE_X26Y131_BO5),
.O6(CLBLL_R_X17Y131_SLICE_X26Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLL_R_X17Y131_SLICE_X26Y131_ALUT (
.I0(1'b1),
.I1(\counter [24]),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y131_SLICE_X26Y131_AO5),
.O6(CLBLL_R_X17Y131_SLICE_X26Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y131_SLICE_X27Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y131_SLICE_X27Y131_DO5),
.O6(CLBLL_R_X17Y131_SLICE_X27Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y131_SLICE_X27Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y131_SLICE_X27Y131_CO5),
.O6(CLBLL_R_X17Y131_SLICE_X27Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y131_SLICE_X27Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y131_SLICE_X27Y131_BO5),
.O6(CLBLL_R_X17Y131_SLICE_X27Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y131_SLICE_X27Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y131_SLICE_X27Y131_AO5),
.O6(CLBLL_R_X17Y131_SLICE_X27Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y132_SLICE_X26Y132_A_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y132_SLICE_X26Y132_A_XOR),
.Q(CLBLL_R_X17Y132_SLICE_X26Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y132_SLICE_X26Y132_B_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y132_SLICE_X26Y132_BO5),
.Q(CLBLL_R_X17Y132_SLICE_X26Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y132_SLICE_X26Y132_C_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y132_SLICE_X26Y132_CO5),
.Q(CLBLL_R_X17Y132_SLICE_X26Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y132_SLICE_X26Y132_D_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y132_SLICE_X26Y132_DO5),
.Q(CLBLL_R_X17Y132_SLICE_X26Y132_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y132_SLICE_X26Y132_CARRY4 (
.CI(\$abc$3569$aiger3568$109 ),
.CO({\$abc$3569$aiger3568$118 , CLBLL_R_X17Y132_SLICE_X26Y132_C_CY, CLBLL_R_X17Y132_SLICE_X26Y132_B_CY, CLBLL_R_X17Y132_SLICE_X26Y132_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1385.O [31], \$auto$alumacc.cc:485:replace_alu$1385.O [30], \$auto$alumacc.cc:485:replace_alu$1385.O [29], CLBLL_R_X17Y132_SLICE_X26Y132_A_XOR}),
.S({CLBLL_R_X17Y132_SLICE_X26Y132_DO6, CLBLL_R_X17Y132_SLICE_X26Y132_CO6, CLBLL_R_X17Y132_SLICE_X26Y132_BO6, CLBLL_R_X17Y132_SLICE_X26Y132_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ff00)
  ) CLBLL_R_X17Y132_SLICE_X26Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_R_X17Y132_SLICE_X26Y132_CQ),
.I3(\$auto$alumacc.cc:485:replace_alu$1385.O [29]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y132_SLICE_X26Y132_DO5),
.O6(CLBLL_R_X17Y132_SLICE_X26Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLL_R_X17Y132_SLICE_X26Y132_CLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1385.O [31]),
.I1(CLBLL_R_X17Y132_SLICE_X26Y132_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y132_SLICE_X26Y132_CO5),
.O6(CLBLL_R_X17Y132_SLICE_X26Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLL_R_X17Y132_SLICE_X26Y132_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X17Y132_SLICE_X26Y132_DQ),
.I2(1'b1),
.I3(\$auto$alumacc.cc:485:replace_alu$1385.O [30]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y132_SLICE_X26Y132_BO5),
.O6(CLBLL_R_X17Y132_SLICE_X26Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLL_R_X17Y132_SLICE_X26Y132_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X17Y132_SLICE_X26Y132_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y132_SLICE_X26Y132_AO5),
.O6(CLBLL_R_X17Y132_SLICE_X26Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y132_SLICE_X27Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y132_SLICE_X27Y132_DO5),
.O6(CLBLL_R_X17Y132_SLICE_X27Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y132_SLICE_X27Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y132_SLICE_X27Y132_CO5),
.O6(CLBLL_R_X17Y132_SLICE_X27Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y132_SLICE_X27Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y132_SLICE_X27Y132_BO5),
.O6(CLBLL_R_X17Y132_SLICE_X27Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y132_SLICE_X27Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y132_SLICE_X27Y132_AO5),
.O6(CLBLL_R_X17Y132_SLICE_X27Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y133_SLICE_X26Y133_A_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y133_SLICE_X26Y133_A_XOR),
.Q(CLBLL_R_X17Y133_SLICE_X26Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y133_SLICE_X26Y133_B_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y133_SLICE_X26Y133_BO5),
.Q(CLBLL_R_X17Y133_SLICE_X26Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y133_SLICE_X26Y133_C_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y133_SLICE_X26Y133_CO5),
.Q(CLBLL_R_X17Y133_SLICE_X26Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y133_SLICE_X26Y133_D_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y133_SLICE_X26Y133_DO5),
.Q(CLBLL_R_X17Y133_SLICE_X26Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y133_SLICE_X26Y133_CARRY4 (
.CI(\$abc$3569$aiger3568$118 ),
.CO({CLBLL_R_X17Y133_SLICE_X26Y133_D_CY, CLBLL_R_X17Y133_SLICE_X26Y133_C_CY, CLBLL_R_X17Y133_SLICE_X26Y133_B_CY, CLBLL_R_X17Y133_SLICE_X26Y133_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1385.O [35], \$auto$alumacc.cc:485:replace_alu$1385.O [34], \$auto$alumacc.cc:485:replace_alu$1385.O [33], CLBLL_R_X17Y133_SLICE_X26Y133_A_XOR}),
.S({CLBLL_R_X17Y133_SLICE_X26Y133_DO6, CLBLL_R_X17Y133_SLICE_X26Y133_CO6, CLBLL_R_X17Y133_SLICE_X26Y133_BO6, CLBLL_R_X17Y133_SLICE_X26Y133_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ff00)
  ) CLBLL_R_X17Y133_SLICE_X26Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_R_X17Y133_SLICE_X26Y133_CQ),
.I3(\$auto$alumacc.cc:485:replace_alu$1385.O [33]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y133_SLICE_X26Y133_DO5),
.O6(CLBLL_R_X17Y133_SLICE_X26Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLL_R_X17Y133_SLICE_X26Y133_CLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1385.O [35]),
.I1(CLBLL_R_X17Y133_SLICE_X26Y133_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y133_SLICE_X26Y133_CO5),
.O6(CLBLL_R_X17Y133_SLICE_X26Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLL_R_X17Y133_SLICE_X26Y133_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X17Y133_SLICE_X26Y133_DQ),
.I2(1'b1),
.I3(\$auto$alumacc.cc:485:replace_alu$1385.O [34]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y133_SLICE_X26Y133_BO5),
.O6(CLBLL_R_X17Y133_SLICE_X26Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLL_R_X17Y133_SLICE_X26Y133_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X17Y133_SLICE_X26Y133_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y133_SLICE_X26Y133_AO5),
.O6(CLBLL_R_X17Y133_SLICE_X26Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y133_SLICE_X27Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y133_SLICE_X27Y133_DO5),
.O6(CLBLL_R_X17Y133_SLICE_X27Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y133_SLICE_X27Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y133_SLICE_X27Y133_CO5),
.O6(CLBLL_R_X17Y133_SLICE_X27Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y133_SLICE_X27Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y133_SLICE_X27Y133_BO5),
.O6(CLBLL_R_X17Y133_SLICE_X27Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y133_SLICE_X27Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y133_SLICE_X27Y133_AO5),
.O6(CLBLL_R_X17Y133_SLICE_X27Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X43Y75_IOB_X1Y76_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O),
.O(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y1_OBUF (
.I(CLBLL_R_X17Y133_SLICE_X26Y133_CQ),
.O(led[7])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y2_OBUF (
.I(CLBLL_R_X17Y133_SLICE_X26Y133_BQ),
.O(led[6])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y121_IOB_X0Y122_IBUF (
.I(sw[3]),
.O(LIOB33_X0Y121_IOB_X0Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y123_IOB_X0Y123_IBUF (
.I(sw[2]),
.O(LIOB33_X0Y123_IOB_X0Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y123_IOB_X0Y124_IBUF (
.I(sw[1]),
.O(LIOB33_X0Y123_IOB_X0Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y125_IOB_X0Y125_IBUF (
.I(sw[0]),
.O(LIOB33_X0Y125_IOB_X0Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y125_IOB_X0Y126_IBUF (
.I(sw[7]),
.O(LIOB33_X0Y125_IOB_X0Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y127_IOB_X0Y127_IBUF (
.I(sw[6]),
.O(LIOB33_X0Y127_IOB_X0Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(sw[5]),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y137_IOB_X0Y137_IBUF (
.I(sw[4]),
.O(LIOB33_X0Y137_IOB_X0Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y51_IOB_X1Y51_OBUF (
.I(CLBLL_R_X17Y133_SLICE_X26Y133_AQ),
.O(led[4])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y51_IOB_X1Y52_OBUF (
.I(CLBLL_R_X17Y132_SLICE_X26Y132_CQ),
.O(led[3])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y55_IOB_X1Y55_OBUF (
.I(CLBLL_R_X17Y132_SLICE_X26Y132_BQ),
.O(led[2])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y57_IOB_X1Y58_OBUF (
.I(CLBLL_R_X17Y132_SLICE_X26Y132_DQ),
.O(led[1])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y61_IOB_X1Y61_OBUF (
.I(CLBLL_R_X17Y132_SLICE_X26Y132_AQ),
.O(led[0])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y75_IOB_X1Y76_IBUF (
.I(clk),
.O(RIOB33_X43Y75_IOB_X1Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_SING_X43Y50_IOB_X1Y50_OBUF (
.I(CLBLL_R_X17Y133_SLICE_X26Y133_DQ),
.O(led[5])
  );
  assign CLBLL_R_X17Y125_SLICE_X26Y125_COUT = \$abc$3569$aiger3568$55 ;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_AQ = \counter [0];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_BQ = \counter [2];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_CQ = \counter [3];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_DQ = \counter [1];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_BMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [1];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_CMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [2];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_DMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [3];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_COUT = \$abc$3569$aiger3568$64 ;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_AQ = \counter [6];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_BQ = \counter [7];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_CQ = \counter [4];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_DQ = \counter [5];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_AMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [4];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_BMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [5];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_CMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [6];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_DMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [7];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_COUT = \$abc$3569$aiger3568$73 ;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_AQ = \counter [10];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_BQ = \counter [11];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_CQ = \counter [8];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_DQ = \counter [9];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_AMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [8];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_BMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [9];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_CMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [10];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_DMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [11];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_COUT = \$abc$3569$aiger3568$82 ;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_AQ = \counter [14];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_BQ = \counter [15];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_CQ = \counter [12];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_DQ = \counter [13];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_AMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [12];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_BMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [13];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_CMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [14];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_DMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [15];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_COUT = \$abc$3569$aiger3568$91 ;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_AQ = \counter [16];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_BQ = \counter [18];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_CQ = \counter [19];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_DQ = \counter [17];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_BMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [17];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_CMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [18];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_DMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [19];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_COUT = \$abc$3569$aiger3568$100 ;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_AQ = \counter [20];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_BQ = \counter [22];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_CQ = \counter [23];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_DQ = \counter [21];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_BMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [21];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_CMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [22];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_DMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [23];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_COUT = \$abc$3569$aiger3568$109 ;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_AQ = \counter [24];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_BQ = \counter [26];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_CQ = \counter [27];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_DQ = \counter [25];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_BMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [25];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_CMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [26];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_DMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [27];
  assign CLBLL_R_X17Y132_SLICE_X26Y132_COUT = \$abc$3569$aiger3568$118 ;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_BMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [29];
  assign CLBLL_R_X17Y132_SLICE_X26Y132_CMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [30];
  assign CLBLL_R_X17Y132_SLICE_X26Y132_DMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [31];
  assign CLBLL_R_X17Y133_SLICE_X26Y133_BMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [33];
  assign CLBLL_R_X17Y133_SLICE_X26Y133_CMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [34];
  assign CLBLL_R_X17Y133_SLICE_X26Y133_DMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [35];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_B_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [1];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_C_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [2];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_D_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [3];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_D_CY = \$abc$3569$aiger3568$55 ;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_A_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [4];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_B_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [5];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_C_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [6];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_D_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [7];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_D_CY = \$abc$3569$aiger3568$64 ;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_A_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [8];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_B_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [9];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_C_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [10];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_D_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [11];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_D_CY = \$abc$3569$aiger3568$73 ;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_A_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [12];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_B_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [13];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_C_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [14];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [15];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D_CY = \$abc$3569$aiger3568$82 ;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_B_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [17];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_C_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [18];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [19];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D_CY = \$abc$3569$aiger3568$91 ;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_B_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [21];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_C_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [22];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_D_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [23];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_D_CY = \$abc$3569$aiger3568$100 ;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_B_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [25];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_C_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [26];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_D_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [27];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_D_CY = \$abc$3569$aiger3568$109 ;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_B_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [29];
  assign CLBLL_R_X17Y132_SLICE_X26Y132_C_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [30];
  assign CLBLL_R_X17Y132_SLICE_X26Y132_D_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [31];
  assign CLBLL_R_X17Y132_SLICE_X26Y132_D_CY = \$abc$3569$aiger3568$118 ;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_B_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [33];
  assign CLBLL_R_X17Y133_SLICE_X26Y133_C_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [34];
  assign CLBLL_R_X17Y133_SLICE_X26Y133_D_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [35];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_A = CLBLL_R_X17Y125_SLICE_X26Y125_AO6;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_B = CLBLL_R_X17Y125_SLICE_X26Y125_BO6;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_C = CLBLL_R_X17Y125_SLICE_X26Y125_CO6;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_D = CLBLL_R_X17Y125_SLICE_X26Y125_DO6;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_A = CLBLL_R_X17Y125_SLICE_X27Y125_AO6;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_B = CLBLL_R_X17Y125_SLICE_X27Y125_BO6;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_C = CLBLL_R_X17Y125_SLICE_X27Y125_CO6;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_D = CLBLL_R_X17Y125_SLICE_X27Y125_DO6;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_A = CLBLL_R_X17Y126_SLICE_X26Y126_AO6;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_B = CLBLL_R_X17Y126_SLICE_X26Y126_BO6;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_C = CLBLL_R_X17Y126_SLICE_X26Y126_CO6;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_D = CLBLL_R_X17Y126_SLICE_X26Y126_DO6;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_A = CLBLL_R_X17Y126_SLICE_X27Y126_AO6;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_B = CLBLL_R_X17Y126_SLICE_X27Y126_BO6;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_C = CLBLL_R_X17Y126_SLICE_X27Y126_CO6;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_D = CLBLL_R_X17Y126_SLICE_X27Y126_DO6;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_A = CLBLL_R_X17Y127_SLICE_X26Y127_AO6;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_B = CLBLL_R_X17Y127_SLICE_X26Y127_BO6;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_C = CLBLL_R_X17Y127_SLICE_X26Y127_CO6;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_D = CLBLL_R_X17Y127_SLICE_X26Y127_DO6;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_A = CLBLL_R_X17Y127_SLICE_X27Y127_AO6;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_B = CLBLL_R_X17Y127_SLICE_X27Y127_BO6;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_C = CLBLL_R_X17Y127_SLICE_X27Y127_CO6;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_D = CLBLL_R_X17Y127_SLICE_X27Y127_DO6;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_A = CLBLL_R_X17Y128_SLICE_X26Y128_AO6;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_B = CLBLL_R_X17Y128_SLICE_X26Y128_BO6;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_C = CLBLL_R_X17Y128_SLICE_X26Y128_CO6;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D = CLBLL_R_X17Y128_SLICE_X26Y128_DO6;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_A = CLBLL_R_X17Y128_SLICE_X27Y128_AO6;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_B = CLBLL_R_X17Y128_SLICE_X27Y128_BO6;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_C = CLBLL_R_X17Y128_SLICE_X27Y128_CO6;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_D = CLBLL_R_X17Y128_SLICE_X27Y128_DO6;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_A = CLBLL_R_X17Y129_SLICE_X26Y129_AO6;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_B = CLBLL_R_X17Y129_SLICE_X26Y129_BO6;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_C = CLBLL_R_X17Y129_SLICE_X26Y129_CO6;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D = CLBLL_R_X17Y129_SLICE_X26Y129_DO6;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_A = CLBLL_R_X17Y129_SLICE_X27Y129_AO6;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_B = CLBLL_R_X17Y129_SLICE_X27Y129_BO6;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_C = CLBLL_R_X17Y129_SLICE_X27Y129_CO6;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_D = CLBLL_R_X17Y129_SLICE_X27Y129_DO6;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_A = CLBLL_R_X17Y130_SLICE_X26Y130_AO6;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_B = CLBLL_R_X17Y130_SLICE_X26Y130_BO6;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_C = CLBLL_R_X17Y130_SLICE_X26Y130_CO6;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_D = CLBLL_R_X17Y130_SLICE_X26Y130_DO6;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_A = CLBLL_R_X17Y130_SLICE_X27Y130_AO6;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_B = CLBLL_R_X17Y130_SLICE_X27Y130_BO6;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_C = CLBLL_R_X17Y130_SLICE_X27Y130_CO6;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_D = CLBLL_R_X17Y130_SLICE_X27Y130_DO6;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_A = CLBLL_R_X17Y131_SLICE_X26Y131_AO6;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_B = CLBLL_R_X17Y131_SLICE_X26Y131_BO6;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_C = CLBLL_R_X17Y131_SLICE_X26Y131_CO6;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_D = CLBLL_R_X17Y131_SLICE_X26Y131_DO6;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_A = CLBLL_R_X17Y131_SLICE_X27Y131_AO6;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_B = CLBLL_R_X17Y131_SLICE_X27Y131_BO6;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_C = CLBLL_R_X17Y131_SLICE_X27Y131_CO6;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_D = CLBLL_R_X17Y131_SLICE_X27Y131_DO6;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_A = CLBLL_R_X17Y132_SLICE_X26Y132_AO6;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_B = CLBLL_R_X17Y132_SLICE_X26Y132_BO6;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_C = CLBLL_R_X17Y132_SLICE_X26Y132_CO6;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_D = CLBLL_R_X17Y132_SLICE_X26Y132_DO6;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_A = CLBLL_R_X17Y132_SLICE_X27Y132_AO6;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_B = CLBLL_R_X17Y132_SLICE_X27Y132_BO6;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_C = CLBLL_R_X17Y132_SLICE_X27Y132_CO6;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_D = CLBLL_R_X17Y132_SLICE_X27Y132_DO6;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_A = CLBLL_R_X17Y133_SLICE_X26Y133_AO6;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_B = CLBLL_R_X17Y133_SLICE_X26Y133_BO6;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_C = CLBLL_R_X17Y133_SLICE_X26Y133_CO6;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_D = CLBLL_R_X17Y133_SLICE_X26Y133_DO6;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_A = CLBLL_R_X17Y133_SLICE_X27Y133_AO6;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_B = CLBLL_R_X17Y133_SLICE_X27Y133_BO6;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_C = CLBLL_R_X17Y133_SLICE_X27Y133_CO6;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_D = CLBLL_R_X17Y133_SLICE_X27Y133_DO6;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_OQ = CLBLL_R_X17Y133_SLICE_X26Y133_BQ;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_TQ = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_OQ = CLBLL_R_X17Y133_SLICE_X26Y133_CQ;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_TQ = 1'b1;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_O = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_O = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_O = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_O = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_OQ = CLBLL_R_X17Y132_SLICE_X26Y132_CQ;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_TQ = 1'b1;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_OQ = CLBLL_R_X17Y133_SLICE_X26Y133_AQ;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_TQ = 1'b1;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_OQ = CLBLL_R_X17Y132_SLICE_X26Y132_BQ;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_TQ = 1'b1;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_OQ = CLBLL_R_X17Y132_SLICE_X26Y132_AQ;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_TQ = 1'b1;
  assign RIOI3_X43Y75_ILOGIC_X1Y76_O = RIOB33_X43Y75_IOB_X1Y76_I;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_OQ = CLBLL_R_X17Y133_SLICE_X26Y133_DQ;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_OQ = CLBLL_R_X17Y132_SLICE_X26Y132_DQ;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_TQ = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_D4 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_B1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_B2 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_B3 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_B4 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_B5 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_B6 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_D5 = 1'b1;
  assign CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_CE = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_D6 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_C1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_C2 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_C3 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_C4 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_C5 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_C6 = 1'b1;
  assign LIOB33_X0Y1_IOB_X0Y1_O = CLBLL_R_X17Y133_SLICE_X26Y133_CQ;
  assign LIOB33_X0Y1_IOB_X0Y2_O = CLBLL_R_X17Y133_SLICE_X26Y133_BQ;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_D1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_D2 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_D3 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_D4 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_D5 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_D6 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_A1 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_A2 = CLBLL_R_X17Y132_SLICE_X26Y132_AQ;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_A3 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_A4 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_A5 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_A6 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_AX = 1'b0;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_B1 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_B2 = CLBLL_R_X17Y132_SLICE_X26Y132_DQ;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_B3 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_B4 = \$auto$alumacc.cc:485:replace_alu$1385.O [30];
  assign CLBLL_R_X17Y132_SLICE_X26Y132_B5 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_B6 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_BX = 1'b0;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_C1 = \$auto$alumacc.cc:485:replace_alu$1385.O [31];
  assign CLBLL_R_X17Y132_SLICE_X26Y132_C2 = CLBLL_R_X17Y132_SLICE_X26Y132_BQ;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_C3 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_C4 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_C5 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_C6 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_CIN = \$abc$3569$aiger3568$109 ;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_CX = 1'b0;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_D1 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_D2 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_D3 = CLBLL_R_X17Y132_SLICE_X26Y132_CQ;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_D4 = \$auto$alumacc.cc:485:replace_alu$1385.O [29];
  assign CLBLL_R_X17Y132_SLICE_X26Y132_D5 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_D6 = 1'b1;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_D = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_DX = 1'b0;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_D1 = CLBLL_R_X17Y132_SLICE_X26Y132_BQ;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_A1 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_A2 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_A3 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_A4 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_A5 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_T1 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_B1 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_B2 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_B3 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_B4 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_B5 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_B6 = 1'b1;
  assign RIOB33_X43Y57_IOB_X1Y58_O = CLBLL_R_X17Y132_SLICE_X26Y132_DQ;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_C1 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_C2 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_C3 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_C4 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_A1 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_A2 = \counter [16];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_A3 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_A4 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_A5 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_A6 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_C5 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_C6 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_AX = 1'b0;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_B1 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_B2 = \counter [17];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_B3 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_B4 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_B5 = \$auto$alumacc.cc:485:replace_alu$1385.O [18];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_B6 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_D1 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_D2 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_BX = 1'b0;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_D3 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_C1 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_C2 = \$auto$alumacc.cc:485:replace_alu$1385.O [19];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_C3 = \counter [18];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_C4 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_C5 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_C6 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_CIN = \$abc$3569$aiger3568$82 ;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_CX = 1'b0;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D1 = \$auto$alumacc.cc:485:replace_alu$1385.O [17];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D2 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D3 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D4 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D5 = \counter [19];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D6 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_DX = 1'b0;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_A1 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_A2 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_A3 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_A4 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_A5 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_A6 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_B1 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_B2 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_B3 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_B4 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_B5 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_B6 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_C1 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_C2 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_C3 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_C4 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_A1 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_A2 = \counter [4];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_A3 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_A4 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_A5 = \$auto$alumacc.cc:485:replace_alu$1385.O [6];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_A6 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_C5 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_C6 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_AX = 1'b0;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_B1 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_B2 = \counter [5];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_B3 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_B4 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_B5 = \$auto$alumacc.cc:485:replace_alu$1385.O [7];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_B6 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_D1 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_D2 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_BX = 1'b0;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_D3 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_C1 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_C2 = \$auto$alumacc.cc:485:replace_alu$1385.O [4];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_C3 = \counter [6];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_C4 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_C5 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_C6 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_CIN = \$abc$3569$aiger3568$55 ;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_CX = 1'b0;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_D1 = \$auto$alumacc.cc:485:replace_alu$1385.O [5];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_D2 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_D3 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_D4 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_D5 = \counter [7];
  assign CLBLL_R_X17Y126_SLICE_X26Y126_D6 = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_D = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_DX = 1'b0;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_A1 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_A2 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_A3 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_A4 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_A5 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_A6 = 1'b1;
  assign RIOB33_X43Y51_IOB_X1Y51_O = CLBLL_R_X17Y133_SLICE_X26Y133_AQ;
  assign RIOB33_X43Y51_IOB_X1Y52_O = CLBLL_R_X17Y132_SLICE_X26Y132_CQ;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_B1 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_B2 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_B3 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_B4 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_B5 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_B6 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_C1 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_C2 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_C3 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_C4 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_C5 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_C6 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_D5 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_D1 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_D2 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_D3 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_D4 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_D5 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_D6 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_D6 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_A1 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_A2 = CLBLL_R_X17Y133_SLICE_X26Y133_AQ;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_A3 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_A4 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_A5 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_A6 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE0 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE1 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_AX = 1'b0;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE0 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_B1 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_B2 = CLBLL_R_X17Y133_SLICE_X26Y133_DQ;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_B3 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_B4 = \$auto$alumacc.cc:485:replace_alu$1385.O [34];
  assign CLBLL_R_X17Y133_SLICE_X26Y133_B5 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_B6 = 1'b1;
  assign RIOB33_SING_X43Y50_IOB_X1Y50_O = CLBLL_R_X17Y133_SLICE_X26Y133_DQ;
  assign RIOI3_X43Y75_ILOGIC_X1Y76_D = RIOB33_X43Y75_IOB_X1Y76_I;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_BX = 1'b0;
  assign CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_I = CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_C1 = \$auto$alumacc.cc:485:replace_alu$1385.O [35];
  assign CLBLL_R_X17Y133_SLICE_X26Y133_C2 = CLBLL_R_X17Y133_SLICE_X26Y133_BQ;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_C3 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_C4 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_C5 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_C6 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_CIN = \$abc$3569$aiger3568$118 ;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_CX = 1'b0;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_D1 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_D2 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_D3 = CLBLL_R_X17Y133_SLICE_X26Y133_CQ;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_D4 = \$auto$alumacc.cc:485:replace_alu$1385.O [33];
  assign CLBLL_R_X17Y133_SLICE_X26Y133_D5 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_D6 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X26Y133_DX = 1'b0;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_A1 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_A2 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_A3 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_A4 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_A5 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_A6 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_B1 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_B2 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_B3 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_B4 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_B5 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_B6 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_D4 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_C1 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_C2 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_C3 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_D5 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_A1 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_A2 = \counter [20];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_A3 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_A4 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_D6 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_A5 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_A6 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_C4 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_AX = 1'b0;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_C5 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_B1 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_B2 = \counter [21];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_B3 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_B4 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_B5 = \$auto$alumacc.cc:485:replace_alu$1385.O [22];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_B6 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_D1 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_BX = 1'b0;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_D2 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_C1 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_C2 = \$auto$alumacc.cc:485:replace_alu$1385.O [23];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_C3 = \counter [22];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_C4 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_C5 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_C6 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_C6 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_CIN = \$abc$3569$aiger3568$91 ;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_CX = 1'b0;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_D1 = \$auto$alumacc.cc:485:replace_alu$1385.O [21];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_D2 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_D3 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_D4 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_D5 = \counter [23];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_D6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_D4 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_DX = 1'b0;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_D5 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_D6 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_A1 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_A2 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_A3 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_A4 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_A5 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_A6 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_B1 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_B2 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_B3 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_B4 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_B5 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_B6 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_D3 = 1'b1;
  assign CLBLL_R_X17Y133_SLICE_X27Y133_D4 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_C1 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_C2 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_C3 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_C4 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_A1 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_A2 = \counter [8];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_A3 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_A4 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_A5 = \$auto$alumacc.cc:485:replace_alu$1385.O [10];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_A6 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_C5 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_C6 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_AX = 1'b0;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_B1 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_B2 = \counter [9];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_B3 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_B4 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_B5 = \$auto$alumacc.cc:485:replace_alu$1385.O [11];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_B6 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_D1 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_D2 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_BX = 1'b0;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_D3 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_C1 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_C2 = \$auto$alumacc.cc:485:replace_alu$1385.O [8];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_C3 = \counter [10];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_C4 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_C5 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_C6 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_CIN = \$abc$3569$aiger3568$64 ;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_D1 = CLBLL_R_X17Y132_SLICE_X26Y132_AQ;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_CX = 1'b0;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_D1 = \$auto$alumacc.cc:485:replace_alu$1385.O [9];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_D2 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_D3 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_D4 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_D5 = \counter [11];
  assign CLBLL_R_X17Y127_SLICE_X26Y127_D6 = 1'b1;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_T1 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X26Y127_DX = 1'b0;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_A1 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_A2 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_A3 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_A4 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_A5 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_A6 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_B1 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_B2 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_B3 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_B4 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_B5 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_B6 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_C1 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_C2 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_C3 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_C4 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_C5 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_C6 = 1'b1;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_D1 = CLBLL_R_X17Y132_SLICE_X26Y132_CQ;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_D1 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_D2 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_D3 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_D4 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_D5 = 1'b1;
  assign CLBLL_R_X17Y127_SLICE_X27Y127_D6 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_D1 = CLBLL_R_X17Y133_SLICE_X26Y133_BQ;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE1 = 1'b1;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_T1 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S0 = 1'b1;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_D1 = CLBLL_R_X17Y133_SLICE_X26Y133_AQ;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S1 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_T1 = 1'b1;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_D = LIOB33_X0Y125_IOB_X0Y126_I;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_T1 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_D1 = CLBLL_R_X17Y133_SLICE_X26Y133_CQ;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_D = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_T1 = 1'b1;
  assign RIOB33_X43Y61_IOB_X1Y61_O = CLBLL_R_X17Y132_SLICE_X26Y132_AQ;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_D1 = CLBLL_R_X17Y132_SLICE_X26Y132_DQ;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_A1 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_A2 = \counter [24];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_A3 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_A4 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_A5 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_T1 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_AX = 1'b0;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_B1 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_B2 = \counter [25];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_B3 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_B4 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_B5 = \$auto$alumacc.cc:485:replace_alu$1385.O [26];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_B6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_BX = 1'b0;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_C1 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_C2 = \$auto$alumacc.cc:485:replace_alu$1385.O [27];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_C3 = \counter [26];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_C4 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_C5 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_C6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_CIN = \$abc$3569$aiger3568$100 ;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_CX = 1'b0;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_D1 = \$auto$alumacc.cc:485:replace_alu$1385.O [25];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_D2 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_D3 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_D4 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_D5 = \counter [27];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_D6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_DX = 1'b0;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_D = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_A1 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_A2 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_A3 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_A4 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_A5 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_A6 = 1'b1;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_D = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_B1 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_B2 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_B3 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_B4 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_B5 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_B6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_C1 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_C2 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_C3 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_C4 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_A1 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_A2 = \counter [12];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_A3 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_A4 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_A5 = \$auto$alumacc.cc:485:replace_alu$1385.O [14];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_A6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_C5 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_C6 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_AX = 1'b0;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_B1 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_B2 = \counter [13];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_B3 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_B4 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_B5 = \$auto$alumacc.cc:485:replace_alu$1385.O [15];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_B6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_D1 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_D2 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_BX = 1'b0;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_D3 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_C1 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_C2 = \$auto$alumacc.cc:485:replace_alu$1385.O [12];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_C3 = \counter [14];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_C4 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_C5 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_C6 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_CIN = \$abc$3569$aiger3568$73 ;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign RIOB33_X43Y55_IOB_X1Y55_O = CLBLL_R_X17Y132_SLICE_X26Y132_BQ;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_CX = 1'b0;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D1 = \$auto$alumacc.cc:485:replace_alu$1385.O [13];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D2 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D3 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D4 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D5 = \counter [15];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D6 = 1'b1;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_D1 = CLBLL_R_X17Y133_SLICE_X26Y133_DQ;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_DX = 1'b0;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_T1 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_A1 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_A2 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_A3 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_A4 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_A5 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_A6 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_B1 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_B2 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_B3 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_B4 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_B5 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_B6 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_C1 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_C2 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_C3 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_C4 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_A1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_A2 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_A3 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_A4 = \counter [0];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_A5 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_A6 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_C5 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_C6 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_AX = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_B1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_B2 = \counter [1];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_B3 = \$auto$alumacc.cc:485:replace_alu$1385.O [2];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_B4 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_D4 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_D5 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_D6 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_B5 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_B6 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_D1 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_D2 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_BX = 1'b0;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_D3 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_C1 = \$auto$alumacc.cc:485:replace_alu$1385.O [3];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_C2 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_C3 = \counter [2];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_C4 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_C5 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_C6 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_D4 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_CX = 1'b0;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_D1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_D2 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_D3 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_D4 = \$auto$alumacc.cc:485:replace_alu$1385.O [1];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_D5 = \counter [3];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_D6 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_D5 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_D6 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_DX = 1'b0;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I0 = RIOB33_X43Y75_IOB_X1Y76_I;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_A1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_A2 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_A3 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_A4 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_A5 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_A6 = 1'b1;
endmodule
