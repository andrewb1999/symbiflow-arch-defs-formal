module top(
  input clk,
  input [7:0] sw,
  output [7:0] led
  );
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A1;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A2;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A3;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A4;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_AO5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_AO6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A_CY;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_A_XOR;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B1;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B2;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B3;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B4;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_BO5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_BO6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B_CY;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_B_XOR;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C1;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C2;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C3;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C4;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_CO5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_CO6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C_CY;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_C_XOR;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D1;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D2;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D3;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D4;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_DO5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_DO6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D_CY;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X26Y125_D_XOR;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A1;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A2;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A3;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A4;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A5Q;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_AMUX;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_AO5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_AO6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_AX;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A_CY;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_A_XOR;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B1;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B2;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B3;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B4;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_BMUX;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_BO5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_BO6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_BQ;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_BX;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B_CY;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_B_XOR;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C1;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C2;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C3;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C4;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_CLK;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_CMUX;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_CO5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_CO6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_COUT;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_CQ;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_CX;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C_CY;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_C_XOR;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D1;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D2;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D3;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D4;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_DMUX;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_DO5;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_DO6;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_DQ;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_DX;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D_CY;
  wire [0:0] CLBLL_R_X17Y125_SLICE_X27Y125_D_XOR;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A1;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A2;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A3;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A4;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_AO5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_AO6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A_CY;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_A_XOR;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B1;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B2;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B3;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B4;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_BO5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_BO6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B_CY;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_B_XOR;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C1;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C2;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C3;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C4;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_CO5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_CO6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C_CY;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_C_XOR;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D1;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D2;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D3;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D4;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_DO5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_DO6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D_CY;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X26Y126_D_XOR;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A1;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A2;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A3;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A4;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_AO5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_AO6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_AQ;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_AX;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A_CY;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_A_XOR;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B1;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B2;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B3;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B4;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_BMUX;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_BO5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_BO6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_BQ;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_BX;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B_CY;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_B_XOR;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C1;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C2;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C3;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C4;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_CIN;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_CLK;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_CMUX;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_CO5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_CO6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_COUT;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_CQ;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_CX;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C_CY;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_C_XOR;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D1;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D2;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D3;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D4;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_DMUX;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_DO5;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_DO6;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_DQ;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_DX;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D_CY;
  wire [0:0] CLBLL_R_X17Y126_SLICE_X27Y126_D_XOR;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S1;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_CE;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_I;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_I;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_O;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y2_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_TQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_TQ;
  wire [0:0] RIOB33_SING_X43Y50_IOB_X1Y50_O;
  wire [0:0] RIOB33_X43Y51_IOB_X1Y51_O;
  wire [0:0] RIOB33_X43Y51_IOB_X1Y52_O;
  wire [0:0] RIOB33_X43Y55_IOB_X1Y55_O;
  wire [0:0] RIOB33_X43Y57_IOB_X1Y58_O;
  wire [0:0] RIOB33_X43Y61_IOB_X1Y61_O;
  wire [0:0] RIOB33_X43Y75_IOB_X1Y76_I;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_D1;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_OQ;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_T1;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_TQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_D1;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_OQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_T1;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_TQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_D1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_OQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_T1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_TQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_D1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_OQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_T1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_TQ;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_D1;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_OQ;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_T1;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_TQ;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_D1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_OQ;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_T1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_TQ;
  wire [0:0] RIOI3_X43Y75_ILOGIC_X1Y76_D;
  wire [0:0] RIOI3_X43Y75_ILOGIC_X1Y76_O;
  wire [0:0] \$abc$3422$aiger3421$27 ;
  wire [7:0] \$auto$alumacc.cc:485:replace_alu$1385.O ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y125_SLICE_X26Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y125_SLICE_X26Y125_DO5),
.O6(CLBLL_R_X17Y125_SLICE_X26Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y125_SLICE_X26Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y125_SLICE_X26Y125_CO5),
.O6(CLBLL_R_X17Y125_SLICE_X26Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y125_SLICE_X26Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y125_SLICE_X26Y125_BO5),
.O6(CLBLL_R_X17Y125_SLICE_X26Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y125_SLICE_X26Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y125_SLICE_X26Y125_AO5),
.O6(CLBLL_R_X17Y125_SLICE_X26Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y125_SLICE_X27Y125_A5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y125_SLICE_X27Y125_AO5),
.Q(CLBLL_R_X17Y125_SLICE_X27Y125_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y125_SLICE_X27Y125_B_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y125_SLICE_X27Y125_BO5),
.Q(CLBLL_R_X17Y125_SLICE_X27Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y125_SLICE_X27Y125_C_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y125_SLICE_X27Y125_CO5),
.Q(CLBLL_R_X17Y125_SLICE_X27Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y125_SLICE_X27Y125_D_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y125_SLICE_X27Y125_DO5),
.Q(CLBLL_R_X17Y125_SLICE_X27Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y125_SLICE_X27Y125_CARRY4 (
.CI(1'b0),
.CO({\$abc$3422$aiger3421$27 , CLBLL_R_X17Y125_SLICE_X27Y125_C_CY, CLBLL_R_X17Y125_SLICE_X27Y125_B_CY, CLBLL_R_X17Y125_SLICE_X27Y125_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({\$auto$alumacc.cc:485:replace_alu$1385.O [3], \$auto$alumacc.cc:485:replace_alu$1385.O [2], \$auto$alumacc.cc:485:replace_alu$1385.O [1], CLBLL_R_X17Y125_SLICE_X27Y125_A_XOR}),
.S({CLBLL_R_X17Y125_SLICE_X27Y125_DO6, CLBLL_R_X17Y125_SLICE_X27Y125_CO6, CLBLL_R_X17Y125_SLICE_X27Y125_BO6, \$auto$alumacc.cc:485:replace_alu$1385.O [0]})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00cccccccc)
  ) CLBLL_R_X17Y125_SLICE_X27Y125_DLUT (
.I0(1'b1),
.I1(\$auto$alumacc.cc:485:replace_alu$1385.O [1]),
.I2(1'b1),
.I3(CLBLL_R_X17Y125_SLICE_X27Y125_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y125_SLICE_X27Y125_DO5),
.O6(CLBLL_R_X17Y125_SLICE_X27Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f0f0f0)
  ) CLBLL_R_X17Y125_SLICE_X27Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(\$auto$alumacc.cc:485:replace_alu$1385.O [3]),
.I3(CLBLL_R_X17Y125_SLICE_X27Y125_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y125_SLICE_X27Y125_CO5),
.O6(CLBLL_R_X17Y125_SLICE_X27Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffff0000)
  ) CLBLL_R_X17Y125_SLICE_X27Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_R_X17Y125_SLICE_X27Y125_DQ),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1385.O [2]),
.I5(1'b1),
.O5(CLBLL_R_X17Y125_SLICE_X27Y125_BO5),
.O6(CLBLL_R_X17Y125_SLICE_X27Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffffff00ff00)
  ) CLBLL_R_X17Y125_SLICE_X27Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(\$auto$alumacc.cc:485:replace_alu$1385.O [0]),
.I4(CLBLL_R_X17Y125_SLICE_X27Y125_A5Q),
.I5(1'b1),
.O5(CLBLL_R_X17Y125_SLICE_X27Y125_AO5),
.O6(\$auto$alumacc.cc:485:replace_alu$1385.O [0])
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y126_SLICE_X26Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y126_SLICE_X26Y126_DO5),
.O6(CLBLL_R_X17Y126_SLICE_X26Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y126_SLICE_X26Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y126_SLICE_X26Y126_CO5),
.O6(CLBLL_R_X17Y126_SLICE_X26Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y126_SLICE_X26Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y126_SLICE_X26Y126_BO5),
.O6(CLBLL_R_X17Y126_SLICE_X26Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y126_SLICE_X26Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y126_SLICE_X26Y126_AO5),
.O6(CLBLL_R_X17Y126_SLICE_X26Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y126_SLICE_X27Y126_A_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y126_SLICE_X27Y126_A_XOR),
.Q(CLBLL_R_X17Y126_SLICE_X27Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y126_SLICE_X27Y126_B_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y126_SLICE_X27Y126_BO5),
.Q(CLBLL_R_X17Y126_SLICE_X27Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y126_SLICE_X27Y126_C_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y126_SLICE_X27Y126_CO5),
.Q(CLBLL_R_X17Y126_SLICE_X27Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y126_SLICE_X27Y126_D_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y126_SLICE_X27Y126_DO5),
.Q(CLBLL_R_X17Y126_SLICE_X27Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y126_SLICE_X27Y126_CARRY4 (
.CI(\$abc$3422$aiger3421$27 ),
.CO({CLBLL_R_X17Y126_SLICE_X27Y126_D_CY, CLBLL_R_X17Y126_SLICE_X27Y126_C_CY, CLBLL_R_X17Y126_SLICE_X27Y126_B_CY, CLBLL_R_X17Y126_SLICE_X27Y126_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1385.O [7], \$auto$alumacc.cc:485:replace_alu$1385.O [6], \$auto$alumacc.cc:485:replace_alu$1385.O [5], CLBLL_R_X17Y126_SLICE_X27Y126_A_XOR}),
.S({CLBLL_R_X17Y126_SLICE_X27Y126_DO6, CLBLL_R_X17Y126_SLICE_X27Y126_CO6, CLBLL_R_X17Y126_SLICE_X27Y126_BO6, CLBLL_R_X17Y126_SLICE_X27Y126_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ff00)
  ) CLBLL_R_X17Y126_SLICE_X27Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_R_X17Y126_SLICE_X27Y126_CQ),
.I3(\$auto$alumacc.cc:485:replace_alu$1385.O [5]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y126_SLICE_X27Y126_DO5),
.O6(CLBLL_R_X17Y126_SLICE_X27Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLL_R_X17Y126_SLICE_X27Y126_CLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1385.O [7]),
.I1(CLBLL_R_X17Y126_SLICE_X27Y126_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y126_SLICE_X27Y126_CO5),
.O6(CLBLL_R_X17Y126_SLICE_X27Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLL_R_X17Y126_SLICE_X27Y126_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X17Y126_SLICE_X27Y126_DQ),
.I2(1'b1),
.I3(\$auto$alumacc.cc:485:replace_alu$1385.O [6]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y126_SLICE_X27Y126_BO5),
.O6(CLBLL_R_X17Y126_SLICE_X27Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLL_R_X17Y126_SLICE_X27Y126_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X17Y126_SLICE_X27Y126_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y126_SLICE_X27Y126_AO5),
.O6(CLBLL_R_X17Y126_SLICE_X27Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X43Y75_IOB_X1Y76_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O),
.O(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y1_OBUF (
.I(CLBLL_R_X17Y126_SLICE_X27Y126_CQ),
.O(led[7])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y2_OBUF (
.I(CLBLL_R_X17Y126_SLICE_X27Y126_BQ),
.O(led[6])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y121_IOB_X0Y122_IBUF (
.I(sw[3]),
.O(LIOB33_X0Y121_IOB_X0Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y123_IOB_X0Y123_IBUF (
.I(sw[2]),
.O(LIOB33_X0Y123_IOB_X0Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y123_IOB_X0Y124_IBUF (
.I(sw[1]),
.O(LIOB33_X0Y123_IOB_X0Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y125_IOB_X0Y125_IBUF (
.I(sw[0]),
.O(LIOB33_X0Y125_IOB_X0Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y125_IOB_X0Y126_IBUF (
.I(sw[7]),
.O(LIOB33_X0Y125_IOB_X0Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y127_IOB_X0Y127_IBUF (
.I(sw[6]),
.O(LIOB33_X0Y127_IOB_X0Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(sw[5]),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y137_IOB_X0Y137_IBUF (
.I(sw[4]),
.O(LIOB33_X0Y137_IOB_X0Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y51_IOB_X1Y51_OBUF (
.I(CLBLL_R_X17Y126_SLICE_X27Y126_AQ),
.O(led[4])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y51_IOB_X1Y52_OBUF (
.I(CLBLL_R_X17Y125_SLICE_X27Y125_CQ),
.O(led[3])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y55_IOB_X1Y55_OBUF (
.I(CLBLL_R_X17Y125_SLICE_X27Y125_BQ),
.O(led[2])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y57_IOB_X1Y58_OBUF (
.I(CLBLL_R_X17Y125_SLICE_X27Y125_DQ),
.O(led[1])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y61_IOB_X1Y61_OBUF (
.I(CLBLL_R_X17Y125_SLICE_X27Y125_A5Q),
.O(led[0])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y75_IOB_X1Y76_IBUF (
.I(clk),
.O(RIOB33_X43Y75_IOB_X1Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_SING_X43Y50_IOB_X1Y50_OBUF (
.I(CLBLL_R_X17Y126_SLICE_X27Y126_DQ),
.O(led[5])
  );
  assign CLBLL_R_X17Y125_SLICE_X27Y125_COUT = \$abc$3422$aiger3421$27 ;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_A = \$auto$alumacc.cc:485:replace_alu$1385.O [0];
  assign CLBLL_R_X17Y125_SLICE_X27Y125_BMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [1];
  assign CLBLL_R_X17Y125_SLICE_X27Y125_CMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [2];
  assign CLBLL_R_X17Y125_SLICE_X27Y125_DMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [3];
  assign CLBLL_R_X17Y126_SLICE_X27Y126_BMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [5];
  assign CLBLL_R_X17Y126_SLICE_X27Y126_CMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [6];
  assign CLBLL_R_X17Y126_SLICE_X27Y126_DMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [7];
  assign CLBLL_R_X17Y125_SLICE_X27Y125_AO6 = \$auto$alumacc.cc:485:replace_alu$1385.O [0];
  assign CLBLL_R_X17Y125_SLICE_X27Y125_B_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [1];
  assign CLBLL_R_X17Y125_SLICE_X27Y125_C_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [2];
  assign CLBLL_R_X17Y125_SLICE_X27Y125_D_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [3];
  assign CLBLL_R_X17Y125_SLICE_X27Y125_D_CY = \$abc$3422$aiger3421$27 ;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_B_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [5];
  assign CLBLL_R_X17Y126_SLICE_X27Y126_C_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [6];
  assign CLBLL_R_X17Y126_SLICE_X27Y126_D_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [7];
  assign CLBLL_R_X17Y125_SLICE_X26Y125_A = CLBLL_R_X17Y125_SLICE_X26Y125_AO6;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_B = CLBLL_R_X17Y125_SLICE_X26Y125_BO6;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_C = CLBLL_R_X17Y125_SLICE_X26Y125_CO6;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_D = CLBLL_R_X17Y125_SLICE_X26Y125_DO6;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_B = CLBLL_R_X17Y125_SLICE_X27Y125_BO6;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_C = CLBLL_R_X17Y125_SLICE_X27Y125_CO6;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_D = CLBLL_R_X17Y125_SLICE_X27Y125_DO6;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_AMUX = CLBLL_R_X17Y125_SLICE_X27Y125_A5Q;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_A = CLBLL_R_X17Y126_SLICE_X26Y126_AO6;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_B = CLBLL_R_X17Y126_SLICE_X26Y126_BO6;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_C = CLBLL_R_X17Y126_SLICE_X26Y126_CO6;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_D = CLBLL_R_X17Y126_SLICE_X26Y126_DO6;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_A = CLBLL_R_X17Y126_SLICE_X27Y126_AO6;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_B = CLBLL_R_X17Y126_SLICE_X27Y126_BO6;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_C = CLBLL_R_X17Y126_SLICE_X27Y126_CO6;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_D = CLBLL_R_X17Y126_SLICE_X27Y126_DO6;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_OQ = CLBLL_R_X17Y126_SLICE_X27Y126_BQ;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_TQ = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_OQ = CLBLL_R_X17Y126_SLICE_X27Y126_CQ;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_TQ = 1'b1;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_O = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_O = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_O = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_O = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_OQ = CLBLL_R_X17Y125_SLICE_X27Y125_CQ;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_TQ = 1'b1;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_OQ = CLBLL_R_X17Y126_SLICE_X27Y126_AQ;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_TQ = 1'b1;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_OQ = CLBLL_R_X17Y125_SLICE_X27Y125_BQ;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_TQ = 1'b1;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_OQ = CLBLL_R_X17Y125_SLICE_X27Y125_A5Q;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_TQ = 1'b1;
  assign RIOI3_X43Y75_ILOGIC_X1Y76_O = RIOB33_X43Y75_IOB_X1Y76_I;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_OQ = CLBLL_R_X17Y126_SLICE_X27Y126_DQ;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_OQ = CLBLL_R_X17Y125_SLICE_X27Y125_DQ;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_TQ = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_AX = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_B1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_B2 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_B3 = CLBLL_R_X17Y125_SLICE_X27Y125_DQ;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_B4 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_B5 = \$auto$alumacc.cc:485:replace_alu$1385.O [2];
  assign CLBLL_R_X17Y125_SLICE_X27Y125_B6 = 1'b1;
  assign CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_CE = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_BX = 1'b0;
  assign LIOB33_X0Y1_IOB_X0Y2_O = CLBLL_R_X17Y126_SLICE_X27Y126_BQ;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_C1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_C2 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_C3 = \$auto$alumacc.cc:485:replace_alu$1385.O [3];
  assign CLBLL_R_X17Y125_SLICE_X27Y125_C4 = CLBLL_R_X17Y125_SLICE_X27Y125_BQ;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_C5 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_C6 = 1'b1;
  assign LIOB33_X0Y1_IOB_X0Y1_O = CLBLL_R_X17Y126_SLICE_X27Y126_CQ;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_CX = 1'b0;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_D1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_D2 = \$auto$alumacc.cc:485:replace_alu$1385.O [1];
  assign CLBLL_R_X17Y125_SLICE_X27Y125_D3 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_D4 = CLBLL_R_X17Y125_SLICE_X27Y125_CQ;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_D5 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_D6 = 1'b1;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_D = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_DX = 1'b0;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_D = LIOB33_X0Y125_IOB_X0Y125_I;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_D1 = CLBLL_R_X17Y125_SLICE_X27Y125_A5Q;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_T1 = 1'b1;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_D = LIOB33_X0Y121_IOB_X0Y122_I;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_D1 = CLBLL_R_X17Y125_SLICE_X27Y125_BQ;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_D1 = CLBLL_R_X17Y125_SLICE_X27Y125_CQ;
  assign RIOB33_X43Y57_IOB_X1Y58_O = CLBLL_R_X17Y125_SLICE_X27Y125_DQ;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_T1 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_D1 = CLBLL_R_X17Y126_SLICE_X27Y126_BQ;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_D1 = CLBLL_R_X17Y126_SLICE_X27Y126_AQ;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_T1 = 1'b1;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_T1 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_D1 = CLBLL_R_X17Y126_SLICE_X27Y126_CQ;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_T1 = 1'b1;
  assign RIOB33_X43Y61_IOB_X1Y61_O = CLBLL_R_X17Y125_SLICE_X27Y125_A5Q;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_A1 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_A2 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_A3 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_A4 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_A5 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_D1 = CLBLL_R_X17Y125_SLICE_X27Y125_DQ;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_B1 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_B2 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_B3 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_B4 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_B5 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_T1 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_C1 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_C2 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_C3 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_C4 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_C5 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_C6 = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_D1 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_D2 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_D3 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_D4 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_D5 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X26Y126_D6 = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_D = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_A1 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_A2 = CLBLL_R_X17Y126_SLICE_X27Y126_AQ;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_A3 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_A4 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_A5 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_A6 = 1'b1;
  assign RIOB33_X43Y51_IOB_X1Y51_O = CLBLL_R_X17Y126_SLICE_X27Y126_AQ;
  assign RIOB33_X43Y51_IOB_X1Y52_O = CLBLL_R_X17Y125_SLICE_X27Y125_CQ;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_AX = 1'b0;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_B1 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_B2 = CLBLL_R_X17Y126_SLICE_X27Y126_DQ;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_B3 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_B4 = \$auto$alumacc.cc:485:replace_alu$1385.O [6];
  assign CLBLL_R_X17Y126_SLICE_X27Y126_B5 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_B6 = 1'b1;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_D = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_D = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_BX = 1'b0;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_C1 = \$auto$alumacc.cc:485:replace_alu$1385.O [7];
  assign CLBLL_R_X17Y126_SLICE_X27Y126_C2 = CLBLL_R_X17Y126_SLICE_X27Y126_BQ;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_C3 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_C4 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_C5 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_C6 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_CIN = \$abc$3422$aiger3421$27 ;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_CX = 1'b0;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_D1 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_D2 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_D3 = CLBLL_R_X17Y126_SLICE_X27Y126_CQ;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_D4 = \$auto$alumacc.cc:485:replace_alu$1385.O [5];
  assign CLBLL_R_X17Y126_SLICE_X27Y126_D5 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_D6 = 1'b1;
  assign CLBLL_R_X17Y126_SLICE_X27Y126_DX = 1'b0;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE0 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE1 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE0 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE1 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S0 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S1 = 1'b1;
  assign RIOB33_X43Y55_IOB_X1Y55_O = CLBLL_R_X17Y125_SLICE_X27Y125_BQ;
  assign RIOB33_SING_X43Y50_IOB_X1Y50_O = CLBLL_R_X17Y126_SLICE_X27Y126_DQ;
  assign RIOI3_X43Y75_ILOGIC_X1Y76_D = RIOB33_X43Y75_IOB_X1Y76_I;
  assign CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_I = CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_D1 = CLBLL_R_X17Y126_SLICE_X27Y126_DQ;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_T1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_A1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_A2 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_A3 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_A4 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_A5 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_A6 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_B1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_B2 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_B3 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_B4 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_B5 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_B6 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_C1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_C2 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_C3 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_C4 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_C5 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_C6 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_D1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_D2 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_D3 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_D4 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_D5 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X26Y125_D6 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I0 = RIOB33_X43Y75_IOB_X1Y76_I;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_A1 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_A2 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_A3 = 1'b1;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_A4 = \$auto$alumacc.cc:485:replace_alu$1385.O [0];
  assign CLBLL_R_X17Y125_SLICE_X27Y125_A5 = CLBLL_R_X17Y125_SLICE_X27Y125_A5Q;
  assign CLBLL_R_X17Y125_SLICE_X27Y125_A6 = 1'b1;
endmodule
