module top(
  input clk,
  input [7:0] sw,
  output [7:0] led
  );
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_XOR;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_A;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_A1;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_A2;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_A3;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_A4;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_A5;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_A6;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_AMUX;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_AO5;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_AO6;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_A_CY;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_A_XOR;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_B;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_B1;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_B2;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_B3;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_B4;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_B5;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_B6;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_BO5;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_BO6;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_B_CY;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_B_XOR;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_C;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_C1;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_C2;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_C3;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_C4;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_C5;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_C6;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_CO5;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_CO6;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_C_CY;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_C_XOR;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_D;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_D1;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_D2;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_D3;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_D4;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_D5;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_D6;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_DO5;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_DO6;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_D_CY;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X18Y120_D_XOR;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_A;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_A1;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_A2;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_A3;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_A4;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_A5;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_A6;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_AO5;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_AO6;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_A_CY;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_A_XOR;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_B;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_B1;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_B2;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_B3;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_B4;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_B5;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_B6;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_BO5;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_BO6;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_B_CY;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_B_XOR;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_C;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_C1;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_C2;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_C3;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_C4;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_C5;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_C6;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_CO5;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_CO6;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_C_CY;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_C_XOR;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_D;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_D1;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_D2;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_D3;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_D4;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_D5;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_D6;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_DO5;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_DO6;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_D_CY;
  wire [0:0] CLBLL_R_X13Y120_SLICE_X19Y120_D_XOR;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S1;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_CE;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_I;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_I;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_O;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y2_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_TQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_TQ;
  wire [0:0] RIOB33_SING_X43Y50_IOB_X1Y50_O;
  wire [0:0] RIOB33_X43Y51_IOB_X1Y51_O;
  wire [0:0] RIOB33_X43Y51_IOB_X1Y52_O;
  wire [0:0] RIOB33_X43Y55_IOB_X1Y55_O;
  wire [0:0] RIOB33_X43Y57_IOB_X1Y58_O;
  wire [0:0] RIOB33_X43Y61_IOB_X1Y61_O;
  wire [0:0] RIOB33_X43Y75_IOB_X1Y76_I;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_D1;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_OQ;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_T1;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_TQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_D1;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_OQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_T1;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_TQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_D1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_OQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_T1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_TQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_D1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_OQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_T1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_TQ;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_D1;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_OQ;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_T1;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_TQ;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_D1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_OQ;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_T1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_TQ;
  wire [0:0] RIOI3_X43Y75_ILOGIC_X1Y76_D;
  wire [0:0] RIOI3_X43Y75_ILOGIC_X1Y76_O;
  wire [5:0] \$techmap1848$abc$1841$lut\led[7].A ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc6ccccc00000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_DLUT (
.I0(LIOB33_X0Y121_IOB_X0Y122_I),
.I1(LIOB33_X0Y127_IOB_X0Y127_I),
.I2(LIOB33_X0Y127_IOB_X0Y128_I),
.I3(\$techmap1848$abc$1841$lut\led[7].A [5]),
.I4(LIOB33_X0Y137_IOB_X0Y137_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h99cc99ccbbff4400)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_CLUT (
.I0(\$techmap1848$abc$1841$lut\led[7].A [5]),
.I1(LIOB33_X0Y137_IOB_X0Y137_I),
.I2(1'b1),
.I3(LIOB33_X0Y121_IOB_X0Y122_I),
.I4(LIOB33_X0Y127_IOB_X0Y128_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f000faaaa5555)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_BLUT (
.I0(\$techmap1848$abc$1841$lut\led[7].A [5]),
.I1(1'b1),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(LIOB33_X0Y123_IOB_X0Y124_I),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_BO5),
.O6(\$techmap1848$abc$1841$lut\led[7].A [5])
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff007f80ff00)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_ALUT (
.I0(LIOB33_X0Y127_IOB_X0Y127_I),
.I1(LIOB33_X0Y127_IOB_X0Y128_I),
.I2(LIOB33_X0Y121_IOB_X0Y122_I),
.I3(LIOB33_X0Y125_IOB_X0Y126_I),
.I4(LIOB33_X0Y137_IOB_X0Y137_I),
.I5(\$techmap1848$abc$1841$lut\led[7].A [5]),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X13Y120_SLICE_X18Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X13Y120_SLICE_X18Y120_DO5),
.O6(CLBLL_R_X13Y120_SLICE_X18Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X13Y120_SLICE_X18Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X13Y120_SLICE_X18Y120_CO5),
.O6(CLBLL_R_X13Y120_SLICE_X18Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X13Y120_SLICE_X18Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X13Y120_SLICE_X18Y120_BO5),
.O6(CLBLL_R_X13Y120_SLICE_X18Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffffcccc3333)
  ) CLBLL_R_X13Y120_SLICE_X18Y120_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y123_IOB_X0Y123_I),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y123_IOB_X0Y124_I),
.I5(1'b1),
.O5(CLBLL_R_X13Y120_SLICE_X18Y120_AO5),
.O6(CLBLL_R_X13Y120_SLICE_X18Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X13Y120_SLICE_X19Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X13Y120_SLICE_X19Y120_DO5),
.O6(CLBLL_R_X13Y120_SLICE_X19Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X13Y120_SLICE_X19Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X13Y120_SLICE_X19Y120_CO5),
.O6(CLBLL_R_X13Y120_SLICE_X19Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X13Y120_SLICE_X19Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X13Y120_SLICE_X19Y120_BO5),
.O6(CLBLL_R_X13Y120_SLICE_X19Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X13Y120_SLICE_X19Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X13Y120_SLICE_X19Y120_AO5),
.O6(CLBLL_R_X13Y120_SLICE_X19Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X43Y75_IOB_X1Y76_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O),
.O(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y1_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.O(led[7])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y2_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X1Y120_DO6),
.O(led[6])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y121_IOB_X0Y122_IBUF (
.I(sw[3]),
.O(LIOB33_X0Y121_IOB_X0Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y123_IOB_X0Y123_IBUF (
.I(sw[2]),
.O(LIOB33_X0Y123_IOB_X0Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y123_IOB_X0Y124_IBUF (
.I(sw[1]),
.O(LIOB33_X0Y123_IOB_X0Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y125_IOB_X0Y125_IBUF (
.I(sw[0]),
.O(LIOB33_X0Y125_IOB_X0Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y125_IOB_X0Y126_IBUF (
.I(sw[7]),
.O(LIOB33_X0Y125_IOB_X0Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y127_IOB_X0Y127_IBUF (
.I(sw[6]),
.O(LIOB33_X0Y127_IOB_X0Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(sw[5]),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y137_IOB_X0Y137_IBUF (
.I(sw[4]),
.O(LIOB33_X0Y137_IOB_X0Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y51_IOB_X1Y51_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X1Y120_CO6),
.O(led[4])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y51_IOB_X1Y52_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X1Y120_BO5),
.O(led[3])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y55_IOB_X1Y55_OBUF (
.I(CLBLL_R_X13Y120_SLICE_X18Y120_AO5),
.O(led[2])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y57_IOB_X1Y58_OBUF (
.I(CLBLL_R_X13Y120_SLICE_X18Y120_AO6),
.O(led[1])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y61_IOB_X1Y61_OBUF (
.I(LIOB33_X0Y125_IOB_X0Y125_I),
.O(led[0])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y75_IOB_X1Y76_IBUF (
.I(clk),
.O(RIOB33_X43Y75_IOB_X1Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_SING_X43Y50_IOB_X1Y50_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X1Y120_CO5),
.O(led[5])
  );
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B = \$techmap1848$abc$1841$lut\led[7].A [5];
  assign CLBLL_L_X2Y120_SLICE_X1Y120_BO6 = \$techmap1848$abc$1841$lut\led[7].A [5];
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_AMUX = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_BMUX = CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_CMUX = CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_DMUX = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_A = CLBLL_R_X13Y120_SLICE_X18Y120_AO6;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_B = CLBLL_R_X13Y120_SLICE_X18Y120_BO6;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_C = CLBLL_R_X13Y120_SLICE_X18Y120_CO6;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_D = CLBLL_R_X13Y120_SLICE_X18Y120_DO6;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_AMUX = CLBLL_R_X13Y120_SLICE_X18Y120_AO5;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_A = CLBLL_R_X13Y120_SLICE_X19Y120_AO6;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_B = CLBLL_R_X13Y120_SLICE_X19Y120_BO6;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_C = CLBLL_R_X13Y120_SLICE_X19Y120_CO6;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_D = CLBLL_R_X13Y120_SLICE_X19Y120_DO6;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_OQ = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_TQ = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_OQ = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_TQ = 1'b1;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_O = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_O = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_O = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_O = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_OQ = CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_TQ = 1'b1;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_OQ = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_TQ = 1'b1;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_OQ = CLBLL_R_X13Y120_SLICE_X18Y120_AO5;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_TQ = 1'b1;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_OQ = LIOB33_X0Y125_IOB_X0Y125_I;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_TQ = 1'b1;
  assign RIOI3_X43Y75_ILOGIC_X1Y76_O = RIOB33_X43Y75_IOB_X1Y76_I;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_OQ = CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_OQ = CLBLL_R_X13Y120_SLICE_X18Y120_AO6;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_TQ = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D6 = 1'b1;
  assign CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_CE = 1'b1;
  assign LIOB33_X0Y1_IOB_X0Y1_O = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign LIOB33_X0Y1_IOB_X0Y2_O = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_D = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_D = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A1 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A2 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A3 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A4 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A5 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A6 = \$techmap1848$abc$1841$lut\led[7].A [5];
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B1 = \$techmap1848$abc$1841$lut\led[7].A [5];
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B4 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B6 = 1'b1;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_D1 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C1 = \$techmap1848$abc$1841$lut\led[7].A [5];
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C2 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C4 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C5 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C6 = 1'b1;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_T1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D1 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D2 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D3 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D4 = \$techmap1848$abc$1841$lut\led[7].A [5];
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D5 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D6 = 1'b1;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_D = LIOB33_X0Y121_IOB_X0Y122_I;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_D1 = CLBLL_R_X13Y120_SLICE_X18Y120_AO5;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_D1 = CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  assign RIOB33_X43Y57_IOB_X1Y58_O = CLBLL_R_X13Y120_SLICE_X18Y120_AO6;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_T1 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_A1 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_A2 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_A3 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_A4 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_A5 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_A6 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_D1 = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_B1 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_B2 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_B3 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_B4 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_B5 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_B6 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_T1 = 1'b1;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_D1 = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_C1 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_C2 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_C3 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_C4 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_C5 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_C6 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_D1 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_T1 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_D1 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_D2 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_D3 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_D4 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_D5 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X18Y120_D6 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_T1 = 1'b1;
  assign RIOB33_X43Y61_IOB_X1Y61_O = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_A1 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_A2 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_A3 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_A4 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_A5 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_A6 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_B1 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_B2 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_B3 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_B4 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_B5 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_B6 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_C1 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_C2 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_C3 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_C4 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_C5 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_D1 = CLBLL_R_X13Y120_SLICE_X18Y120_AO6;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_D1 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_D2 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_D3 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_D4 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_D5 = 1'b1;
  assign CLBLL_R_X13Y120_SLICE_X19Y120_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_T1 = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_D = LIOB33_X0Y127_IOB_X0Y127_I;
  assign RIOB33_X43Y51_IOB_X1Y52_O = CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  assign RIOB33_X43Y51_IOB_X1Y51_O = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_D = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_D = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE0 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE1 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE0 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE1 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S0 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S1 = 1'b1;
  assign RIOB33_X43Y55_IOB_X1Y55_O = CLBLL_R_X13Y120_SLICE_X18Y120_AO5;
  assign RIOB33_SING_X43Y50_IOB_X1Y50_O = CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  assign RIOI3_X43Y75_ILOGIC_X1Y76_D = RIOB33_X43Y75_IOB_X1Y76_I;
  assign CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_I = CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_D1 = CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_T1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B6 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I0 = RIOB33_X43Y75_IOB_X1Y76_I;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C6 = 1'b1;
endmodule
