module top(
  input clk,
  input [7:0] sw,
  output [7:0] led
  );
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_A;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_A1;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_A2;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_A3;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_A4;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_A5;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_A6;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_AMUX;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_AO5;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_AO6;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_A_CY;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_A_XOR;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_B;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_B1;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_B2;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_B3;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_B4;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_B5;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_B5Q;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_B6;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_BMUX;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_BO5;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_BO6;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_BQ;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_BX;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_B_CY;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_B_XOR;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_C;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_C1;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_C2;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_C3;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_C4;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_C5;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_C5Q;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_C6;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_CLK;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_CMUX;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_CO5;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_CO6;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_CQ;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_CX;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_C_CY;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_C_XOR;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_D;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_D1;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_D2;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_D3;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_D4;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_D5;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_D5Q;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_D6;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_DMUX;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_DO5;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_DO6;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_DQ;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_DX;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_D_CY;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X18Y135_D_XOR;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_A;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_A1;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_A2;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_A3;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_A4;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_A5;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_A6;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_AMUX;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_AO5;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_AO6;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_A_CY;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_A_XOR;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_B;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_B1;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_B2;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_B3;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_B4;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_B5;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_B6;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_BMUX;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_BO5;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_BO6;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_B_CY;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_B_XOR;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_C;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_C1;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_C2;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_C3;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_C4;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_C5;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_C5Q;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_C6;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_CLK;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_CMUX;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_CO5;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_CO6;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_CQ;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_CX;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_C_CY;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_C_XOR;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_D;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_D1;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_D2;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_D3;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_D4;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_D5;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_D6;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_DMUX;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_DO5;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_DO6;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_D_CY;
  wire [0:0] CLBLL_R_X13Y135_SLICE_X19Y135_D_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_AO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_AO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_BO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_BO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_CO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_CO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_DO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_DO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_AMUX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_AO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_AO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_BMUX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_BO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_BO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C5Q;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CLK;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CMUX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CQ;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D5Q;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_DMUX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_DO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_DO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_DQ;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_DX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D_XOR;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A1;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A2;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A3;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A4;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_AMUX;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_AO5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_AO6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A_CY;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_A_XOR;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B1;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B2;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B3;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B4;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_BMUX;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_BO5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_BO6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_BQ;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_BX;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B_CY;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_B_XOR;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C1;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C2;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C3;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C4;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C5Q;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_CLK;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_CMUX;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_CO5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_CO6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_CQ;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_CX;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C_CY;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_C_XOR;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D1;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D2;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D3;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D4;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D5Q;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_DMUX;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_DO5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_DO6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_DQ;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_DX;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D_CY;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X26Y128_D_XOR;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A1;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A2;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A3;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A4;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_AO5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_AO6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A_CY;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_A_XOR;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B1;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B2;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B3;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B4;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_BO5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_BO6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B_CY;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_B_XOR;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C1;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C2;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C3;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C4;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_CO5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_CO6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C_CY;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_C_XOR;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D1;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D2;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D3;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D4;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_DO5;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_DO6;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D_CY;
  wire [0:0] CLBLL_R_X17Y128_SLICE_X27Y128_D_XOR;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A1;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A2;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A3;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A4;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_AMUX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_AO5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_AO6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A_CY;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_A_XOR;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B1;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B2;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B3;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B4;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_BMUX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_BO5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_BO6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_BQ;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_BX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B_CY;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_B_XOR;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C1;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C2;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C3;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C4;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C5Q;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_CLK;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_CMUX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_CO5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_CO6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_CQ;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_CX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C_CY;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_C_XOR;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D1;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D2;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D3;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D4;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D5Q;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_DMUX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_DO5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_DO6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_DX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D_CY;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X26Y129_D_XOR;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A1;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A2;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A3;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A4;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_AMUX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_AO5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_AO6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_AQ;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_AX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A_CY;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_A_XOR;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B1;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B2;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B3;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B4;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_BMUX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_BO5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_BO6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B_CY;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_B_XOR;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C1;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C2;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C3;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C4;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C5Q;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_CLK;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_CMUX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_CO5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_CO6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_CX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C_CY;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_C_XOR;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D1;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D2;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D3;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D4;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_DMUX;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_DO5;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_DO6;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D_CY;
  wire [0:0] CLBLL_R_X17Y129_SLICE_X27Y129_D_XOR;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A1;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A2;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A3;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A4;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_AMUX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_AO5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_AO6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_AQ;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_AX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A_CY;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_A_XOR;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B1;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B2;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B3;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B4;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_BMUX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_BO5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_BO6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_BQ;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_BX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B_CY;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_B_XOR;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C1;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C2;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C3;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C4;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C5Q;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_CLK;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_CMUX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_CO5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_CO6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_CQ;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_CX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C_CY;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_C_XOR;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D1;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D2;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D3;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D4;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_DMUX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_DO5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_DO6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D_CY;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X26Y130_D_XOR;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A1;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A2;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A3;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A4;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_AMUX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_AO5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_AO6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A_CY;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_A_XOR;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B1;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B2;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B3;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B4;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_BMUX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_BO5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_BO6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B_CY;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_B_XOR;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C1;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C2;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C3;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C4;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C5Q;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_CLK;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_CMUX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_CO5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_CO6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_CQ;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_CX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C_CY;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_C_XOR;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D1;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D2;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D3;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D4;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_DMUX;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_DO5;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_DO6;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D_CY;
  wire [0:0] CLBLL_R_X17Y130_SLICE_X27Y130_D_XOR;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A1;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A2;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A3;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A4;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_AMUX;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_AO5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_AO6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A_CY;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_A_XOR;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B1;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B2;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B3;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B4;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_BO5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_BO6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B_CY;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_B_XOR;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C1;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C2;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C3;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C4;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_CO5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_CO6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C_CY;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_C_XOR;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D1;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D2;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D3;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D4;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_DO5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_DO6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D_CY;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X26Y131_D_XOR;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A1;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A2;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A3;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A4;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_AMUX;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_AO5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_AO6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A_CY;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_A_XOR;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B1;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B2;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B3;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B4;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_BMUX;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_BO5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_BO6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B_CY;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_B_XOR;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C1;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C2;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C3;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C4;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C5Q;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_CLK;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_CMUX;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_CO5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_CO6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_CQ;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_CX;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C_CY;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_C_XOR;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D1;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D2;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D3;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D4;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D5Q;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_DMUX;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_DO5;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_DO6;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_DX;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D_CY;
  wire [0:0] CLBLL_R_X17Y131_SLICE_X27Y131_D_XOR;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A1;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A2;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A3;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A4;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_AO5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_AO6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A_CY;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_A_XOR;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B1;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B2;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B3;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B4;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_BO5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_BO6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B_CY;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_B_XOR;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C1;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C2;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C3;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C4;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_CO5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_CO6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C_CY;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_C_XOR;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D1;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D2;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D3;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D4;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_DO5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_DO6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D_CY;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X26Y132_D_XOR;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A1;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A2;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A3;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A4;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_AMUX;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_AO5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_AO6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_AQ;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A_CY;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_A_XOR;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B1;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B2;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B3;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B4;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_BMUX;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_BO5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_BO6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_BQ;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B_CY;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_B_XOR;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C1;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C2;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C3;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C4;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C5Q;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_CLK;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_CMUX;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_CO5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_CO6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_CQ;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_CX;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C_CY;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_C_XOR;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D1;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D2;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D3;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D4;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_DMUX;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_DO5;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_DO6;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D_CY;
  wire [0:0] CLBLL_R_X17Y132_SLICE_X27Y132_D_XOR;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S1;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_CE;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_I;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_I;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_O;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y2_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_TQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_TQ;
  wire [0:0] RIOB33_SING_X43Y50_IOB_X1Y50_O;
  wire [0:0] RIOB33_X43Y51_IOB_X1Y51_O;
  wire [0:0] RIOB33_X43Y51_IOB_X1Y52_O;
  wire [0:0] RIOB33_X43Y55_IOB_X1Y55_O;
  wire [0:0] RIOB33_X43Y57_IOB_X1Y58_O;
  wire [0:0] RIOB33_X43Y61_IOB_X1Y61_O;
  wire [0:0] RIOB33_X43Y75_IOB_X1Y76_I;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_D1;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_OQ;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_T1;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_TQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_D1;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_OQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_T1;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_TQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_D1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_OQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_T1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_TQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_D1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_OQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_T1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_TQ;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_D1;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_OQ;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_T1;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_TQ;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_D1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_OQ;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_T1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_TQ;
  wire [0:0] RIOI3_X43Y75_ILOGIC_X1Y76_D;
  wire [0:0] RIOI3_X43Y75_ILOGIC_X1Y76_O;
  wire [0:0] \$auto$alumacc.cc:485:replace_alu$1415.X ;
  wire [35:0] \$auto$alumacc.cc:485:replace_alu$1415.Y ;
  wire [5:0] \$techmap2792$abc$2783$lut$aiger2782$78.A ;
  wire [3:0] \$techmap2797$abc$2783$lut$aiger2782$68.A ;
  wire [1:0] \$techmap2798$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[6].A ;
  wire [2:0] \$techmap2807$abc$2783$lut$aiger2782$226.A ;
  wire [5:0] \$techmap2810$abc$2783$lut$aiger2782$176.A ;
  wire [3:0] \$techmap2812$abc$2783$lut$aiger2782$119.A ;
  wire [5:0] \$techmap2813$abc$2783$lut$aiger2782$231.A ;
  wire [3:0] \$techmap2819$abc$2783$lut$aiger2782$187.A ;
  wire [4:0] \$techmap2820$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[30].A ;
  wire [5:0] \$techmap2822$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[29].A ;
  wire [1:0] \$techmap2829$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[23].A ;
  wire [3:0] \$techmap2834$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[20].A ;
  wire [2:0] \$techmap2839$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[16].A ;
  wire [2:0] \$techmap2843$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[13].A ;
  wire [27:0] \counter ;


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1505CLBLL_R_X13Y135_SLICE_X18Y135_B5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [5]),
.Q(\counter [5]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1507CLBLL_R_X13Y135_SLICE_X18Y135_C5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X13Y135_SLICE_X18Y135_CO5),
.Q(\counter [7]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1506CLBLL_R_X13Y135_SLICE_X18Y135_D5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [6]),
.Q(\counter [6]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1501CLBLL_R_X13Y135_SLICE_X18Y135_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X13Y135_SLICE_X18Y135_BO5),
.Q(\counter [1]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1503CLBLL_R_X13Y135_SLICE_X18Y135_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [3]),
.Q(\counter [3]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1502CLBLL_R_X13Y135_SLICE_X18Y135_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X13Y135_SLICE_X18Y135_DO5),
.Q(\counter [2]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ffff0000)
  ) CLBLL_R_X13Y135_SLICE_X18Y135_DLUT (
.I0(1'b1),
.I1(\counter [3]),
.I2(1'b1),
.I3(\$techmap2792$abc$2783$lut$aiger2782$78.A [5]),
.I4(\$auto$alumacc.cc:485:replace_alu$1415.Y [2]),
.I5(1'b1),
.O5(CLBLL_R_X13Y135_SLICE_X18Y135_DO5),
.O6(\$techmap2797$abc$2783$lut$aiger2782$68.A [3])
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88008800ffff0000)
  ) CLBLL_R_X13Y135_SLICE_X18Y135_CLUT (
.I0(\counter [2]),
.I1(\counter [0]),
.I2(1'b1),
.I3(\counter [1]),
.I4(\$auto$alumacc.cc:485:replace_alu$1415.Y [7]),
.I5(1'b1),
.O5(CLBLL_R_X13Y135_SLICE_X18Y135_CO5),
.O6(\$techmap2792$abc$2783$lut$aiger2782$78.A [5])
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff03333cccc)
  ) CLBLL_R_X13Y135_SLICE_X18Y135_BLUT (
.I0(1'b1),
.I1(\counter [1]),
.I2(\counter [7]),
.I3(\$techmap2798$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[6].A [1]),
.I4(\counter [0]),
.I5(1'b1),
.O5(CLBLL_R_X13Y135_SLICE_X18Y135_BO5),
.O6(\$auto$alumacc.cc:485:replace_alu$1415.Y [7])
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_R_X13Y135_SLICE_X18Y135_ALUT (
.I0(\counter [7]),
.I1(\counter [6]),
.I2(\counter [3]),
.I3(\counter [4]),
.I4(\counter [5]),
.I5(\$techmap2792$abc$2783$lut$aiger2782$78.A [5]),
.O5(CLBLL_R_X13Y135_SLICE_X18Y135_AO5),
.O6(CLBLL_R_X13Y135_SLICE_X18Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1504CLBLL_R_X13Y135_SLICE_X19Y135_C5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X13Y135_SLICE_X19Y135_CO5),
.Q(\counter [4]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1500CLBLL_R_X13Y135_SLICE_X19Y135_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.X [0]),
.Q(\counter [0]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0ff000f0f0f0f)
  ) CLBLL_R_X13Y135_SLICE_X19Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(\counter [0]),
.I3(\counter [2]),
.I4(\counter [1]),
.I5(1'b1),
.O5(\$auto$alumacc.cc:485:replace_alu$1415.X [0]),
.O6(\$auto$alumacc.cc:485:replace_alu$1415.Y [2])
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h66666666ff00ff00)
  ) CLBLL_R_X13Y135_SLICE_X19Y135_CLUT (
.I0(\$techmap2792$abc$2783$lut$aiger2782$78.A [5]),
.I1(\counter [3]),
.I2(1'b1),
.I3(\$auto$alumacc.cc:485:replace_alu$1415.Y [4]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X13Y135_SLICE_X19Y135_CO5),
.O6(\$auto$alumacc.cc:485:replace_alu$1415.Y [3])
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5af0f05fa0ff00)
  ) CLBLL_R_X13Y135_SLICE_X19Y135_BLUT (
.I0(\$techmap2797$abc$2783$lut$aiger2782$68.A [3]),
.I1(1'b1),
.I2(\counter [5]),
.I3(\counter [6]),
.I4(\counter [4]),
.I5(1'b1),
.O5(\$auto$alumacc.cc:485:replace_alu$1415.Y [6]),
.O6(\$auto$alumacc.cc:485:replace_alu$1415.Y [5])
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha00000005a5a5a5a)
  ) CLBLL_R_X13Y135_SLICE_X19Y135_ALUT (
.I0(\$techmap2797$abc$2783$lut$aiger2782$68.A [3]),
.I1(1'b1),
.I2(\counter [4]),
.I3(\counter [5]),
.I4(\counter [6]),
.I5(1'b1),
.O5(\$auto$alumacc.cc:485:replace_alu$1415.Y [4]),
.O6(\$techmap2798$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[6].A [1])
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y120_SLICE_X26Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X26Y120_DO5),
.O6(CLBLL_R_X17Y120_SLICE_X26Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y120_SLICE_X26Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X26Y120_CO5),
.O6(CLBLL_R_X17Y120_SLICE_X26Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y120_SLICE_X26Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X26Y120_BO5),
.O6(CLBLL_R_X17Y120_SLICE_X26Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y120_SLICE_X26Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X26Y120_AO5),
.O6(CLBLL_R_X17Y120_SLICE_X26Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_C5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y120_SLICE_X27Y120_CO5),
.Q(CLBLL_R_X17Y120_SLICE_X27Y120_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_D5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y120_SLICE_X27Y120_DO5),
.Q(CLBLL_R_X17Y120_SLICE_X27Y120_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_C_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [33]),
.Q(CLBLL_R_X17Y120_SLICE_X27Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_D_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [35]),
.Q(CLBLL_R_X17Y120_SLICE_X27Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_DLUT (
.I0(1'b1),
.I1(\$auto$alumacc.cc:485:replace_alu$1415.Y [34]),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X27Y120_DO5),
.O6(CLBLL_R_X17Y120_SLICE_X27Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaaaaaa)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_CLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1415.Y [32]),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X27Y120_CO5),
.O6(CLBLL_R_X17Y120_SLICE_X27Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5af0f0f06ccccccc)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_BLUT (
.I0(CLBLL_R_X17Y120_SLICE_X27Y120_CQ),
.I1(CLBLL_R_X17Y120_SLICE_X27Y120_DQ),
.I2(CLBLL_R_X17Y120_SLICE_X27Y120_D5Q),
.I3(CLBLL_R_X17Y130_SLICE_X27Y130_BO6),
.I4(CLBLL_R_X17Y120_SLICE_X27Y120_C5Q),
.I5(1'b1),
.O5(\$auto$alumacc.cc:485:replace_alu$1415.Y [35]),
.O6(\$auto$alumacc.cc:485:replace_alu$1415.Y [34])
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cccccc00ffff00)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X17Y120_SLICE_X27Y120_CQ),
.I2(1'b1),
.I3(CLBLL_R_X17Y130_SLICE_X27Y130_BO6),
.I4(CLBLL_R_X17Y120_SLICE_X27Y120_C5Q),
.I5(1'b1),
.O5(\$auto$alumacc.cc:485:replace_alu$1415.Y [32]),
.O6(\$auto$alumacc.cc:485:replace_alu$1415.Y [33])
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y128_SLICE_X26Y128_C5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y128_SLICE_X26Y128_CO5),
.Q(CLBLL_R_X17Y128_SLICE_X26Y128_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1526CLBLL_R_X17Y128_SLICE_X26Y128_D5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y128_SLICE_X26Y128_DO5),
.Q(\counter [26]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y128_SLICE_X26Y128_B_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [28]),
.Q(CLBLL_R_X17Y128_SLICE_X26Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1527CLBLL_R_X17Y128_SLICE_X26Y128_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [27]),
.Q(\counter [27]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y128_SLICE_X26Y128_D_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y129_SLICE_X27Y129_DO6),
.Q(CLBLL_R_X17Y128_SLICE_X26Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h80808080ffff0000)
  ) CLBLL_R_X17Y128_SLICE_X26Y128_DLUT (
.I0(CLBLL_R_X17Y128_SLICE_X26Y128_BQ),
.I1(CLBLL_R_X17Y128_SLICE_X26Y128_C5Q),
.I2(CLBLL_R_X17Y128_SLICE_X26Y128_DQ),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1415.Y [26]),
.I5(1'b1),
.O5(CLBLL_R_X17Y128_SLICE_X26Y128_DO5),
.O6(\$techmap2807$abc$2783$lut$aiger2782$226.A [1])
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aaff00f0f0f0f0)
  ) CLBLL_R_X17Y128_SLICE_X26Y128_CLUT (
.I0(\$techmap2822$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[29].A [5]),
.I1(1'b1),
.I2(CLBLL_R_X17Y128_SLICE_X26Y128_AO6),
.I3(\counter [26]),
.I4(\counter [25]),
.I5(1'b1),
.O5(CLBLL_R_X17Y128_SLICE_X26Y128_CO5),
.O6(\$auto$alumacc.cc:485:replace_alu$1415.Y [26])
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f00078f078f0)
  ) CLBLL_R_X17Y128_SLICE_X26Y128_BLUT (
.I0(\$techmap2822$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[29].A [5]),
.I1(\counter [25]),
.I2(\counter [27]),
.I3(\counter [26]),
.I4(1'b1),
.I5(1'b1),
.O5(\$auto$alumacc.cc:485:replace_alu$1415.Y [27]),
.O6(\$techmap2807$abc$2783$lut$aiger2782$226.A [2])
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6aaaaaaaaaaaaaaa)
  ) CLBLL_R_X17Y128_SLICE_X26Y128_ALUT (
.I0(CLBLL_R_X17Y128_SLICE_X26Y128_C5Q),
.I1(CLBLL_R_X17Y128_SLICE_X26Y128_DQ),
.I2(CLBLL_R_X17Y128_SLICE_X26Y128_BQ),
.I3(\counter [25]),
.I4(\$techmap2807$abc$2783$lut$aiger2782$226.A [2]),
.I5(\$techmap2822$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[29].A [5]),
.O5(CLBLL_R_X17Y128_SLICE_X26Y128_AO5),
.O6(CLBLL_R_X17Y128_SLICE_X26Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y128_SLICE_X27Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y128_SLICE_X27Y128_DO5),
.O6(CLBLL_R_X17Y128_SLICE_X27Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y128_SLICE_X27Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y128_SLICE_X27Y128_CO5),
.O6(CLBLL_R_X17Y128_SLICE_X27Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y128_SLICE_X27Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y128_SLICE_X27Y128_BO5),
.O6(CLBLL_R_X17Y128_SLICE_X27Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y128_SLICE_X27Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y128_SLICE_X27Y128_AO5),
.O6(CLBLL_R_X17Y128_SLICE_X27Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y129_SLICE_X26Y129_C5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y129_SLICE_X26Y129_CO5),
.Q(CLBLL_R_X17Y129_SLICE_X26Y129_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1520CLBLL_R_X17Y129_SLICE_X26Y129_D5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [20]),
.Q(\counter [20]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1517CLBLL_R_X17Y129_SLICE_X26Y129_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [17]),
.Q(\counter [17]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1521CLBLL_R_X17Y129_SLICE_X26Y129_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [21]),
.Q(\counter [21]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000000000000000)
  ) CLBLL_R_X17Y129_SLICE_X26Y129_DLUT (
.I0(\counter [17]),
.I1(1'b1),
.I2(CLBLL_R_X13Y135_SLICE_X18Y135_AO6),
.I3(\$techmap2819$abc$2783$lut$aiger2782$187.A [3]),
.I4(\counter [16]),
.I5(1'b1),
.O5(CLBLL_R_X17Y129_SLICE_X26Y129_DO5),
.O6(\$techmap2834$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[20].A [3])
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f0f0f0f0)
  ) CLBLL_R_X17Y129_SLICE_X26Y129_CLUT (
.I0(1'b1),
.I1(\counter [16]),
.I2(\$auto$alumacc.cc:485:replace_alu$1415.Y [31]),
.I3(\counter [17]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y129_SLICE_X26Y129_CO5),
.O6(\$techmap2810$abc$2783$lut$aiger2782$176.A [5])
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fffa0005af05af0)
  ) CLBLL_R_X17Y129_SLICE_X26Y129_BLUT (
.I0(\$techmap2810$abc$2783$lut$aiger2782$176.A [4]),
.I1(1'b1),
.I2(\counter [20]),
.I3(\$techmap2834$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[20].A [3]),
.I4(\counter [21]),
.I5(1'b1),
.O5(\$auto$alumacc.cc:485:replace_alu$1415.Y [20]),
.O6(\$auto$alumacc.cc:485:replace_alu$1415.Y [21])
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00000007fff8000)
  ) CLBLL_R_X17Y129_SLICE_X26Y129_ALUT (
.I0(\counter [25]),
.I1(\$techmap2820$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[30].A [4]),
.I2(\$techmap2807$abc$2783$lut$aiger2782$226.A [1]),
.I3(\$techmap2807$abc$2783$lut$aiger2782$226.A [2]),
.I4(CLBLL_R_X17Y129_SLICE_X26Y129_C5Q),
.I5(1'b1),
.O5(\$auto$alumacc.cc:485:replace_alu$1415.Y [31]),
.O6(\$techmap2813$abc$2783$lut$aiger2782$231.A [2])
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1525CLBLL_R_X17Y129_SLICE_X27Y129_C5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [25]),
.Q(\counter [25]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1515CLBLL_R_X17Y129_SLICE_X27Y129_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [15]),
.Q(\counter [15]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ccccccc00000000)
  ) CLBLL_R_X17Y129_SLICE_X27Y129_DLUT (
.I0(CLBLL_R_X17Y128_SLICE_X26Y128_BQ),
.I1(CLBLL_R_X17Y128_SLICE_X26Y128_DQ),
.I2(\$techmap2807$abc$2783$lut$aiger2782$226.A [2]),
.I3(\counter [25]),
.I4(\$techmap2822$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[29].A [5]),
.I5(1'b1),
.O5(CLBLL_R_X17Y129_SLICE_X27Y129_DO5),
.O6(CLBLL_R_X17Y129_SLICE_X27Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000000000000)
  ) CLBLL_R_X17Y129_SLICE_X27Y129_CLUT (
.I0(\$techmap2812$abc$2783$lut$aiger2782$119.A [3]),
.I1(\counter [15]),
.I2(1'b1),
.I3(\counter [14]),
.I4(\$techmap2812$abc$2783$lut$aiger2782$119.A [2]),
.I5(1'b1),
.O5(CLBLL_R_X17Y129_SLICE_X27Y129_CO5),
.O6(\$techmap2819$abc$2783$lut$aiger2782$187.A [3])
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080000088000000)
  ) CLBLL_R_X17Y129_SLICE_X27Y129_BLUT (
.I0(\counter [24]),
.I1(CLBLL_R_X17Y130_SLICE_X27Y130_AO6),
.I2(\$techmap2813$abc$2783$lut$aiger2782$231.A [5]),
.I3(\$techmap2819$abc$2783$lut$aiger2782$187.A [3]),
.I4(CLBLL_R_X13Y135_SLICE_X18Y135_AO6),
.I5(1'b1),
.O5(\$techmap2820$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[30].A [4]),
.O6(\$techmap2822$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[29].A [5])
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ff880055aa55aa)
  ) CLBLL_R_X17Y129_SLICE_X27Y129_ALUT (
.I0(\$techmap2822$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[29].A [5]),
.I1(\$techmap2807$abc$2783$lut$aiger2782$226.A [2]),
.I2(1'b1),
.I3(\counter [25]),
.I4(CLBLL_R_X17Y128_SLICE_X26Y128_BQ),
.I5(1'b1),
.O5(\$auto$alumacc.cc:485:replace_alu$1415.Y [25]),
.O6(\$auto$alumacc.cc:485:replace_alu$1415.Y [28])
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1516CLBLL_R_X17Y130_SLICE_X26Y130_C5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [16]),
.Q(\counter [16]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1514CLBLL_R_X17Y130_SLICE_X26Y130_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [14]),
.Q(\counter [14]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1512CLBLL_R_X17Y130_SLICE_X26Y130_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [12]),
.Q(\counter [12]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1513CLBLL_R_X17Y130_SLICE_X26Y130_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y130_SLICE_X26Y130_CO6),
.Q(\counter [13]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f80ff00aaaa0000)
  ) CLBLL_R_X17Y130_SLICE_X26Y130_DLUT (
.I0(CLBLL_R_X13Y135_SLICE_X18Y135_AO6),
.I1(\counter [14]),
.I2(\$techmap2812$abc$2783$lut$aiger2782$119.A [2]),
.I3(\counter [15]),
.I4(\$techmap2812$abc$2783$lut$aiger2782$119.A [3]),
.I5(1'b1),
.O5(\$techmap2843$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[13].A [2]),
.O6(\$auto$alumacc.cc:485:replace_alu$1415.Y [15])
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ccc3ccc00000000)
  ) CLBLL_R_X17Y130_SLICE_X26Y130_CLUT (
.I0(1'b1),
.I1(\counter [13]),
.I2(\$techmap2843$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[13].A [2]),
.I3(\counter [12]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y130_SLICE_X26Y130_CO5),
.O6(CLBLL_R_X17Y130_SLICE_X26Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff0cccc0000)
  ) CLBLL_R_X17Y130_SLICE_X26Y130_BLUT (
.I0(1'b1),
.I1(\counter [13]),
.I2(\counter [18]),
.I3(\$techmap2834$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[20].A [3]),
.I4(\counter [12]),
.I5(1'b1),
.O5(\$techmap2812$abc$2783$lut$aiger2782$119.A [2]),
.O6(\$auto$alumacc.cc:485:replace_alu$1415.Y [18])
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c6c6c6c5a5a5a5a)
  ) CLBLL_R_X17Y130_SLICE_X26Y130_ALUT (
.I0(\$techmap2839$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[16].A [2]),
.I1(\counter [17]),
.I2(\counter [16]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(\$auto$alumacc.cc:485:replace_alu$1415.Y [16]),
.O6(\$auto$alumacc.cc:485:replace_alu$1415.Y [17])
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1519CLBLL_R_X17Y130_SLICE_X27Y130_C5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y130_SLICE_X27Y130_CO5),
.Q(\counter [19]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1518CLBLL_R_X17Y130_SLICE_X27Y130_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [18]),
.Q(\counter [18]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_R_X17Y130_SLICE_X27Y130_DLUT (
.I0(\counter [21]),
.I1(\counter [20]),
.I2(\$techmap2810$abc$2783$lut$aiger2782$176.A [5]),
.I3(\$techmap2810$abc$2783$lut$aiger2782$176.A [4]),
.I4(CLBLL_R_X13Y135_SLICE_X18Y135_AO6),
.I5(\$techmap2813$abc$2783$lut$aiger2782$231.A [5]),
.O5(CLBLL_R_X17Y130_SLICE_X27Y130_DO5),
.O6(CLBLL_R_X17Y130_SLICE_X27Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa005aaa5aaa)
  ) CLBLL_R_X17Y130_SLICE_X27Y130_CLUT (
.I0(\counter [19]),
.I1(1'b1),
.I2(\$techmap2834$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[20].A [3]),
.I3(\counter [18]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y130_SLICE_X27Y130_CO5),
.O6(\$techmap2810$abc$2783$lut$aiger2782$176.A [4])
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_R_X17Y130_SLICE_X27Y130_BLUT (
.I0(\counter [25]),
.I1(CLBLL_R_X13Y135_SLICE_X18Y135_AO6),
.I2(\$techmap2813$abc$2783$lut$aiger2782$231.A [2]),
.I3(CLBLL_R_X17Y130_SLICE_X27Y130_AO6),
.I4(\counter [24]),
.I5(\$techmap2813$abc$2783$lut$aiger2782$231.A [5]),
.O5(CLBLL_R_X17Y130_SLICE_X27Y130_BO5),
.O6(CLBLL_R_X17Y130_SLICE_X27Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_R_X17Y130_SLICE_X27Y130_ALUT (
.I0(\counter [22]),
.I1(\$techmap2810$abc$2783$lut$aiger2782$176.A [4]),
.I2(\counter [23]),
.I3(\counter [21]),
.I4(\counter [20]),
.I5(\$techmap2810$abc$2783$lut$aiger2782$176.A [5]),
.O5(CLBLL_R_X17Y130_SLICE_X27Y130_AO5),
.O6(CLBLL_R_X17Y130_SLICE_X27Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y131_SLICE_X26Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y131_SLICE_X26Y131_DO5),
.O6(CLBLL_R_X17Y131_SLICE_X26Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y131_SLICE_X26Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y131_SLICE_X26Y131_CO5),
.O6(CLBLL_R_X17Y131_SLICE_X26Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y131_SLICE_X26Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y131_SLICE_X26Y131_BO5),
.O6(CLBLL_R_X17Y131_SLICE_X26Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaa33cccccc)
  ) CLBLL_R_X17Y131_SLICE_X26Y131_ALUT (
.I0(\counter [12]),
.I1(\counter [14]),
.I2(1'b1),
.I3(\$techmap2812$abc$2783$lut$aiger2782$119.A [2]),
.I4(\$techmap2843$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[13].A [2]),
.I5(1'b1),
.O5(\$auto$alumacc.cc:485:replace_alu$1415.Y [14]),
.O6(\$auto$alumacc.cc:485:replace_alu$1415.Y [12])
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1523CLBLL_R_X17Y131_SLICE_X27Y131_C5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y131_SLICE_X27Y131_CO5),
.Q(\counter [23]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1522CLBLL_R_X17Y131_SLICE_X27Y131_D5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [22]),
.Q(\counter [22]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1524CLBLL_R_X17Y131_SLICE_X27Y131_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$auto$alumacc.cc:485:replace_alu$1415.Y [24]),
.Q(\counter [24]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000000000000)
  ) CLBLL_R_X17Y131_SLICE_X27Y131_DLUT (
.I0(\counter [14]),
.I1(\counter [15]),
.I2(1'b1),
.I3(\$techmap2812$abc$2783$lut$aiger2782$119.A [2]),
.I4(\$techmap2812$abc$2783$lut$aiger2782$119.A [3]),
.I5(1'b1),
.O5(CLBLL_R_X17Y131_SLICE_X27Y131_DO5),
.O6(\$techmap2813$abc$2783$lut$aiger2782$231.A [5])
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0ff00ff00)
  ) CLBLL_R_X17Y131_SLICE_X27Y131_CLUT (
.I0(\$techmap2813$abc$2783$lut$aiger2782$231.A [5]),
.I1(1'b1),
.I2(CLBLL_R_X13Y135_SLICE_X18Y135_AO6),
.I3(\$auto$alumacc.cc:485:replace_alu$1415.Y [23]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y131_SLICE_X27Y131_CO5),
.O6(\$techmap2839$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[16].A [2])
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000000066666666)
  ) CLBLL_R_X17Y131_SLICE_X27Y131_BLUT (
.I0(\counter [22]),
.I1(CLBLL_R_X17Y130_SLICE_X27Y130_DO6),
.I2(CLBLL_R_X17Y130_SLICE_X27Y130_AO6),
.I3(\$techmap2813$abc$2783$lut$aiger2782$231.A [5]),
.I4(CLBLL_R_X13Y135_SLICE_X18Y135_AO6),
.I5(1'b1),
.O5(\$auto$alumacc.cc:485:replace_alu$1415.Y [22]),
.O6(\$techmap2829$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[23].A [1])
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaa54445444)
  ) CLBLL_R_X17Y131_SLICE_X27Y131_ALUT (
.I0(\$techmap2829$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[23].A [1]),
.I1(\counter [23]),
.I2(\counter [22]),
.I3(CLBLL_R_X17Y130_SLICE_X27Y130_DO6),
.I4(\counter [24]),
.I5(1'b1),
.O5(\$auto$alumacc.cc:485:replace_alu$1415.Y [23]),
.O6(\$auto$alumacc.cc:485:replace_alu$1415.Y [24])
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y132_SLICE_X26Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y132_SLICE_X26Y132_DO5),
.O6(CLBLL_R_X17Y132_SLICE_X26Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y132_SLICE_X26Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y132_SLICE_X26Y132_CO5),
.O6(CLBLL_R_X17Y132_SLICE_X26Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y132_SLICE_X26Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y132_SLICE_X26Y132_BO5),
.O6(CLBLL_R_X17Y132_SLICE_X26Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y132_SLICE_X26Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y132_SLICE_X26Y132_AO5),
.O6(CLBLL_R_X17Y132_SLICE_X26Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1508CLBLL_R_X17Y132_SLICE_X27Y132_C5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y132_SLICE_X27Y132_CO5),
.Q(\counter [8]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1509CLBLL_R_X17Y132_SLICE_X27Y132_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y132_SLICE_X27Y132_AO6),
.Q(\counter [9]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1510CLBLL_R_X17Y132_SLICE_X27Y132_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y132_SLICE_X27Y132_BO5),
.Q(\counter [10]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1511CLBLL_R_X17Y132_SLICE_X27Y132_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y132_SLICE_X27Y132_DO6),
.Q(\counter [11]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h78f0f0f000000000)
  ) CLBLL_R_X17Y132_SLICE_X27Y132_DLUT (
.I0(CLBLL_R_X13Y135_SLICE_X18Y135_AO6),
.I1(\counter [8]),
.I2(\counter [11]),
.I3(\counter [9]),
.I4(\counter [10]),
.I5(1'b1),
.O5(CLBLL_R_X17Y132_SLICE_X27Y132_DO5),
.O6(CLBLL_R_X17Y132_SLICE_X27Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLL_R_X17Y132_SLICE_X27Y132_CLUT (
.I0(1'b1),
.I1(CLBLL_R_X17Y132_SLICE_X27Y132_BO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y132_SLICE_X27Y132_CO5),
.O6(CLBLL_R_X17Y132_SLICE_X27Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaa66cccccc)
  ) CLBLL_R_X17Y132_SLICE_X27Y132_BLUT (
.I0(CLBLL_R_X13Y135_SLICE_X18Y135_AO6),
.I1(\counter [10]),
.I2(1'b1),
.I3(\counter [9]),
.I4(\counter [8]),
.I5(1'b1),
.O5(CLBLL_R_X17Y132_SLICE_X27Y132_BO5),
.O6(CLBLL_R_X17Y132_SLICE_X27Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cccccc80008000)
  ) CLBLL_R_X17Y132_SLICE_X27Y132_ALUT (
.I0(\counter [10]),
.I1(\counter [9]),
.I2(\counter [11]),
.I3(\counter [8]),
.I4(CLBLL_R_X13Y135_SLICE_X18Y135_AO6),
.I5(1'b1),
.O5(\$techmap2812$abc$2783$lut$aiger2782$119.A [3]),
.O6(CLBLL_R_X17Y132_SLICE_X27Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X43Y75_IOB_X1Y76_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O),
.O(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y1_OBUF (
.I(CLBLL_R_X17Y120_SLICE_X27Y120_DQ),
.O(led[7])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y2_OBUF (
.I(CLBLL_R_X17Y120_SLICE_X27Y120_D5Q),
.O(led[6])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y121_IOB_X0Y122_IBUF (
.I(sw[3]),
.O(LIOB33_X0Y121_IOB_X0Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y123_IOB_X0Y123_IBUF (
.I(sw[2]),
.O(LIOB33_X0Y123_IOB_X0Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y123_IOB_X0Y124_IBUF (
.I(sw[1]),
.O(LIOB33_X0Y123_IOB_X0Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y125_IOB_X0Y125_IBUF (
.I(sw[0]),
.O(LIOB33_X0Y125_IOB_X0Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y125_IOB_X0Y126_IBUF (
.I(sw[7]),
.O(LIOB33_X0Y125_IOB_X0Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y127_IOB_X0Y127_IBUF (
.I(sw[6]),
.O(LIOB33_X0Y127_IOB_X0Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(sw[5]),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y137_IOB_X0Y137_IBUF (
.I(sw[4]),
.O(LIOB33_X0Y137_IOB_X0Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y51_IOB_X1Y51_OBUF (
.I(CLBLL_R_X17Y120_SLICE_X27Y120_C5Q),
.O(led[4])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y51_IOB_X1Y52_OBUF (
.I(CLBLL_R_X17Y129_SLICE_X26Y129_C5Q),
.O(led[3])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y55_IOB_X1Y55_OBUF (
.I(CLBLL_R_X17Y128_SLICE_X26Y128_C5Q),
.O(led[2])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y57_IOB_X1Y58_OBUF (
.I(CLBLL_R_X17Y128_SLICE_X26Y128_DQ),
.O(led[1])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y61_IOB_X1Y61_OBUF (
.I(CLBLL_R_X17Y128_SLICE_X26Y128_BQ),
.O(led[0])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y75_IOB_X1Y76_IBUF (
.I(clk),
.O(RIOB33_X43Y75_IOB_X1Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_SING_X43Y50_IOB_X1Y50_OBUF (
.I(CLBLL_R_X17Y120_SLICE_X27Y120_CQ),
.O(led[5])
  );
  assign CLBLL_R_X13Y135_SLICE_X18Y135_BQ = \counter [1];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_CQ = \counter [3];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_DQ = \counter [2];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_B = \$auto$alumacc.cc:485:replace_alu$1415.Y [7];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_C = \$techmap2792$abc$2783$lut$aiger2782$78.A [5];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_D = \$techmap2797$abc$2783$lut$aiger2782$68.A [3];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_BMUX = \counter [5];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_CMUX = \counter [7];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_DMUX = \counter [6];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_CQ = \counter [0];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_A = \$techmap2798$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[6].A [1];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_B = \$auto$alumacc.cc:485:replace_alu$1415.Y [5];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_C = \$auto$alumacc.cc:485:replace_alu$1415.Y [3];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_D = \$auto$alumacc.cc:485:replace_alu$1415.Y [2];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_AMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [4];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_BMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [6];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_CMUX = \counter [4];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_DMUX = \$auto$alumacc.cc:485:replace_alu$1415.X [0];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A = \$auto$alumacc.cc:485:replace_alu$1415.Y [33];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B = \$auto$alumacc.cc:485:replace_alu$1415.Y [34];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_AMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [32];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_BMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [35];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_CQ = \counter [27];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_B = \$techmap2807$abc$2783$lut$aiger2782$226.A [2];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_C = \$auto$alumacc.cc:485:replace_alu$1415.Y [26];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D = \$techmap2807$abc$2783$lut$aiger2782$226.A [1];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_BMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [27];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_DMUX = \counter [26];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_BQ = \counter [17];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_CQ = \counter [21];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_A = \$techmap2813$abc$2783$lut$aiger2782$231.A [2];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_B = \$auto$alumacc.cc:485:replace_alu$1415.Y [21];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_C = \$techmap2810$abc$2783$lut$aiger2782$176.A [5];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D = \$techmap2834$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[20].A [3];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_AMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [31];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_BMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [20];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_DMUX = \counter [20];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_AQ = \counter [15];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_A = \$auto$alumacc.cc:485:replace_alu$1415.Y [28];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_B = \$techmap2822$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[29].A [5];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_C = \$techmap2819$abc$2783$lut$aiger2782$187.A [3];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_AMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [25];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_BMUX = \$techmap2820$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[30].A [4];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_CMUX = \counter [25];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_AQ = \counter [14];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_BQ = \counter [12];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_CQ = \counter [13];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_A = \$auto$alumacc.cc:485:replace_alu$1415.Y [17];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_B = \$auto$alumacc.cc:485:replace_alu$1415.Y [18];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_D = \$auto$alumacc.cc:485:replace_alu$1415.Y [15];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_AMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [16];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_BMUX = \$techmap2812$abc$2783$lut$aiger2782$119.A [2];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_CMUX = \counter [16];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_DMUX = \$techmap2843$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[13].A [2];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_CQ = \counter [18];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_C = \$techmap2810$abc$2783$lut$aiger2782$176.A [4];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_CMUX = \counter [19];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_A = \$auto$alumacc.cc:485:replace_alu$1415.Y [12];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_AMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [14];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_CQ = \counter [24];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_A = \$auto$alumacc.cc:485:replace_alu$1415.Y [24];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_B = \$techmap2829$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[23].A [1];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_C = \$techmap2839$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[16].A [2];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_D = \$techmap2813$abc$2783$lut$aiger2782$231.A [5];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_AMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [23];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_BMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [22];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_CMUX = \counter [23];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_DMUX = \counter [22];
  assign CLBLL_R_X17Y132_SLICE_X27Y132_AQ = \counter [9];
  assign CLBLL_R_X17Y132_SLICE_X27Y132_BQ = \counter [10];
  assign CLBLL_R_X17Y132_SLICE_X27Y132_CQ = \counter [11];
  assign CLBLL_R_X17Y132_SLICE_X27Y132_AMUX = \$techmap2812$abc$2783$lut$aiger2782$119.A [3];
  assign CLBLL_R_X17Y132_SLICE_X27Y132_CMUX = \counter [8];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_DO6 = \$techmap2797$abc$2783$lut$aiger2782$68.A [3];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_CO6 = \$techmap2792$abc$2783$lut$aiger2782$78.A [5];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_BO6 = \$auto$alumacc.cc:485:replace_alu$1415.Y [7];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_B5Q = \counter [5];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_C5Q = \counter [7];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_D5Q = \counter [6];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_DO6 = \$auto$alumacc.cc:485:replace_alu$1415.Y [2];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_DO5 = \$auto$alumacc.cc:485:replace_alu$1415.X [0];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_CO6 = \$auto$alumacc.cc:485:replace_alu$1415.Y [3];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_BO6 = \$auto$alumacc.cc:485:replace_alu$1415.Y [5];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_BO5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [6];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_AO6 = \$techmap2798$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[6].A [1];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_AO5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [4];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_C5Q = \counter [4];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_BO6 = \$auto$alumacc.cc:485:replace_alu$1415.Y [34];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_BO5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [35];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_AO6 = \$auto$alumacc.cc:485:replace_alu$1415.Y [33];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_AO5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [32];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_DO6 = \$techmap2807$abc$2783$lut$aiger2782$226.A [1];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_CO6 = \$auto$alumacc.cc:485:replace_alu$1415.Y [26];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_BO6 = \$techmap2807$abc$2783$lut$aiger2782$226.A [2];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_BO5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [27];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D5Q = \counter [26];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_DO6 = \$techmap2834$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[20].A [3];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_CO6 = \$techmap2810$abc$2783$lut$aiger2782$176.A [5];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_BO6 = \$auto$alumacc.cc:485:replace_alu$1415.Y [21];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_BO5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [20];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_AO6 = \$techmap2813$abc$2783$lut$aiger2782$231.A [2];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_AO5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [31];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D5Q = \counter [20];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_CO6 = \$techmap2819$abc$2783$lut$aiger2782$187.A [3];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_BO6 = \$techmap2822$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[29].A [5];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_BO5 = \$techmap2820$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[30].A [4];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_AO6 = \$auto$alumacc.cc:485:replace_alu$1415.Y [28];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_AO5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [25];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_C5Q = \counter [25];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_DO6 = \$auto$alumacc.cc:485:replace_alu$1415.Y [15];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_DO5 = \$techmap2843$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[13].A [2];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_BO6 = \$auto$alumacc.cc:485:replace_alu$1415.Y [18];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_BO5 = \$techmap2812$abc$2783$lut$aiger2782$119.A [2];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_AO6 = \$auto$alumacc.cc:485:replace_alu$1415.Y [17];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_AO5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [16];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_C5Q = \counter [16];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_CO6 = \$techmap2810$abc$2783$lut$aiger2782$176.A [4];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_C5Q = \counter [19];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_AO6 = \$auto$alumacc.cc:485:replace_alu$1415.Y [12];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_AO5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [14];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_DO6 = \$techmap2813$abc$2783$lut$aiger2782$231.A [5];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_CO6 = \$techmap2839$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[16].A [2];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_BO6 = \$techmap2829$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[23].A [1];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_BO5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [22];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_AO6 = \$auto$alumacc.cc:485:replace_alu$1415.Y [24];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_AO5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [23];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_C5Q = \counter [23];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_D5Q = \counter [22];
  assign CLBLL_R_X17Y132_SLICE_X27Y132_AO5 = \$techmap2812$abc$2783$lut$aiger2782$119.A [3];
  assign CLBLL_R_X17Y132_SLICE_X27Y132_C5Q = \counter [8];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_A = CLBLL_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLL_R_X13Y135_SLICE_X18Y135_AMUX = CLBLL_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A = CLBLL_R_X17Y120_SLICE_X26Y120_AO6;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B = CLBLL_R_X17Y120_SLICE_X26Y120_BO6;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C = CLBLL_R_X17Y120_SLICE_X26Y120_CO6;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D = CLBLL_R_X17Y120_SLICE_X26Y120_DO6;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C = CLBLL_R_X17Y120_SLICE_X27Y120_CO6;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D = CLBLL_R_X17Y120_SLICE_X27Y120_DO6;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_CMUX = CLBLL_R_X17Y120_SLICE_X27Y120_C5Q;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_DMUX = CLBLL_R_X17Y120_SLICE_X27Y120_D5Q;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_A = CLBLL_R_X17Y128_SLICE_X26Y128_AO6;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_AMUX = CLBLL_R_X17Y128_SLICE_X26Y128_AO6;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_CMUX = CLBLL_R_X17Y128_SLICE_X26Y128_C5Q;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_A = CLBLL_R_X17Y128_SLICE_X27Y128_AO6;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_B = CLBLL_R_X17Y128_SLICE_X27Y128_BO6;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_C = CLBLL_R_X17Y128_SLICE_X27Y128_CO6;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_D = CLBLL_R_X17Y128_SLICE_X27Y128_DO6;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_CMUX = CLBLL_R_X17Y129_SLICE_X26Y129_C5Q;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_D = CLBLL_R_X17Y129_SLICE_X27Y129_DO6;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_DMUX = CLBLL_R_X17Y129_SLICE_X27Y129_DO6;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_C = CLBLL_R_X17Y130_SLICE_X26Y130_CO6;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_A = CLBLL_R_X17Y130_SLICE_X27Y130_AO6;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_B = CLBLL_R_X17Y130_SLICE_X27Y130_BO6;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_D = CLBLL_R_X17Y130_SLICE_X27Y130_DO6;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_AMUX = CLBLL_R_X17Y130_SLICE_X27Y130_AO6;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_BMUX = CLBLL_R_X17Y130_SLICE_X27Y130_BO6;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_DMUX = CLBLL_R_X17Y130_SLICE_X27Y130_DO6;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_B = CLBLL_R_X17Y131_SLICE_X26Y131_BO6;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_C = CLBLL_R_X17Y131_SLICE_X26Y131_CO6;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_D = CLBLL_R_X17Y131_SLICE_X26Y131_DO6;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_A = CLBLL_R_X17Y132_SLICE_X26Y132_AO6;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_B = CLBLL_R_X17Y132_SLICE_X26Y132_BO6;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_C = CLBLL_R_X17Y132_SLICE_X26Y132_CO6;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_D = CLBLL_R_X17Y132_SLICE_X26Y132_DO6;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_A = CLBLL_R_X17Y132_SLICE_X27Y132_AO6;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_B = CLBLL_R_X17Y132_SLICE_X27Y132_BO6;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_C = CLBLL_R_X17Y132_SLICE_X27Y132_CO6;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_D = CLBLL_R_X17Y132_SLICE_X27Y132_DO6;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_BMUX = CLBLL_R_X17Y132_SLICE_X27Y132_BO6;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_DMUX = CLBLL_R_X17Y132_SLICE_X27Y132_DO6;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_OQ = CLBLL_R_X17Y120_SLICE_X27Y120_D5Q;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_TQ = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_OQ = CLBLL_R_X17Y120_SLICE_X27Y120_DQ;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_TQ = 1'b1;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_O = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_O = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_O = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_O = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_OQ = CLBLL_R_X17Y129_SLICE_X26Y129_C5Q;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_TQ = 1'b1;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_OQ = CLBLL_R_X17Y120_SLICE_X27Y120_C5Q;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_TQ = 1'b1;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_OQ = CLBLL_R_X17Y128_SLICE_X26Y128_C5Q;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_TQ = 1'b1;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_OQ = CLBLL_R_X17Y128_SLICE_X26Y128_BQ;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_TQ = 1'b1;
  assign RIOI3_X43Y75_ILOGIC_X1Y76_O = RIOB33_X43Y75_IOB_X1Y76_I;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_OQ = CLBLL_R_X17Y120_SLICE_X27Y120_CQ;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_OQ = CLBLL_R_X17Y128_SLICE_X26Y128_DQ;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_TQ = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_D4 = \counter [9];
  assign CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_CE = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_D5 = \counter [10];
  assign CLBLL_R_X17Y132_SLICE_X27Y132_D6 = 1'b1;
  assign LIOB33_X0Y1_IOB_X0Y1_O = CLBLL_R_X17Y120_SLICE_X27Y120_DQ;
  assign LIOB33_X0Y1_IOB_X0Y2_O = CLBLL_R_X17Y120_SLICE_X27Y120_D5Q;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_B6 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_A1 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_A2 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_A3 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_C1 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_A4 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_A5 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_A6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_C2 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_B1 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_B2 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_B3 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_C3 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_B4 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_B5 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_B6 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_C1 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_C2 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_C3 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_C4 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_C5 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_C6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_C6 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_D1 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_D2 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_D3 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_D4 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_D5 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X26Y132_D6 = 1'b1;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_D = LIOB33_X0Y121_IOB_X0Y122_I;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_D1 = CLBLL_R_X17Y128_SLICE_X26Y128_C5Q;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_A1 = \counter [10];
  assign CLBLL_R_X17Y132_SLICE_X27Y132_A2 = \counter [9];
  assign CLBLL_R_X17Y132_SLICE_X27Y132_A3 = \counter [11];
  assign CLBLL_R_X17Y132_SLICE_X27Y132_A4 = \counter [8];
  assign CLBLL_R_X17Y132_SLICE_X27Y132_A5 = CLBLL_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_T1 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_B1 = CLBLL_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_B2 = \counter [10];
  assign CLBLL_R_X17Y132_SLICE_X27Y132_B3 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_B4 = \counter [9];
  assign CLBLL_R_X17Y132_SLICE_X27Y132_B5 = \counter [8];
  assign CLBLL_R_X17Y132_SLICE_X27Y132_B6 = 1'b1;
  assign RIOB33_X43Y57_IOB_X1Y58_O = CLBLL_R_X17Y128_SLICE_X26Y128_DQ;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_C1 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_C2 = CLBLL_R_X17Y132_SLICE_X27Y132_BO6;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_C3 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_C4 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_A1 = \counter [25];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_A2 = \$techmap2820$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[30].A [4];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_A3 = \$techmap2807$abc$2783$lut$aiger2782$226.A [1];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_A4 = \$techmap2807$abc$2783$lut$aiger2782$226.A [2];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_A5 = CLBLL_R_X17Y129_SLICE_X26Y129_C5Q;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_A6 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_C5 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_C6 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_B1 = \$techmap2810$abc$2783$lut$aiger2782$176.A [4];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_B2 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_B3 = \counter [20];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_B4 = \$techmap2834$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[20].A [3];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_B5 = \counter [21];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_B6 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_CX = CLBLL_R_X17Y132_SLICE_X27Y132_DO6;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_D1 = CLBLL_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_BX = \$auto$alumacc.cc:485:replace_alu$1415.Y [17];
  assign CLBLL_R_X17Y132_SLICE_X27Y132_D2 = \counter [8];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_C1 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_C2 = \counter [16];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_C3 = \$auto$alumacc.cc:485:replace_alu$1415.Y [31];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_C4 = \counter [17];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_C5 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_C6 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_CX = \$auto$alumacc.cc:485:replace_alu$1415.Y [21];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D1 = \counter [17];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D2 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D3 = CLBLL_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D4 = \$techmap2819$abc$2783$lut$aiger2782$187.A [3];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D5 = \counter [16];
  assign CLBLL_R_X17Y129_SLICE_X26Y129_D6 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X26Y129_DX = \$auto$alumacc.cc:485:replace_alu$1415.Y [20];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_A1 = \$techmap2822$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[29].A [5];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_A2 = \$techmap2807$abc$2783$lut$aiger2782$226.A [2];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_A3 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_A4 = \counter [25];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_A5 = CLBLL_R_X17Y128_SLICE_X26Y128_BQ;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_A6 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_AX = \$auto$alumacc.cc:485:replace_alu$1415.Y [15];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_B1 = \counter [24];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_B2 = CLBLL_R_X17Y130_SLICE_X27Y130_AO6;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_B3 = \$techmap2813$abc$2783$lut$aiger2782$231.A [5];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_B4 = \$techmap2819$abc$2783$lut$aiger2782$187.A [3];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_B5 = CLBLL_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_B6 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_C1 = \$techmap2812$abc$2783$lut$aiger2782$119.A [3];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_C2 = \counter [15];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_C3 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_C4 = \counter [14];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_C5 = \$techmap2812$abc$2783$lut$aiger2782$119.A [2];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_C6 = 1'b1;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_CX = \$auto$alumacc.cc:485:replace_alu$1415.Y [25];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_D1 = CLBLL_R_X17Y128_SLICE_X26Y128_BQ;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_D2 = CLBLL_R_X17Y128_SLICE_X26Y128_DQ;
  assign CLBLL_R_X17Y129_SLICE_X27Y129_D3 = \$techmap2807$abc$2783$lut$aiger2782$226.A [2];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_D4 = \counter [25];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_D5 = \$techmap2822$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[29].A [5];
  assign CLBLL_R_X17Y129_SLICE_X27Y129_D6 = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_D = LIOB33_X0Y127_IOB_X0Y127_I;
  assign RIOB33_X43Y51_IOB_X1Y52_O = CLBLL_R_X17Y129_SLICE_X26Y129_C5Q;
  assign RIOB33_X43Y51_IOB_X1Y51_O = CLBLL_R_X17Y120_SLICE_X27Y120_C5Q;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE0 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE1 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE0 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE1 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S0 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S1 = 1'b1;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_T1 = 1'b1;
  assign RIOB33_SING_X43Y50_IOB_X1Y50_O = CLBLL_R_X17Y120_SLICE_X27Y120_CQ;
  assign RIOI3_X43Y75_ILOGIC_X1Y76_D = RIOB33_X43Y75_IOB_X1Y76_I;
  assign CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_I = CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A2 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B2 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C2 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C6 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_A1 = \$techmap2839$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[16].A [2];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_A2 = \counter [17];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_A3 = \counter [16];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_A4 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_A5 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_A6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D2 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D6 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_AX = \$auto$alumacc.cc:485:replace_alu$1415.Y [14];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_B1 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_B2 = \counter [13];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_B3 = \counter [18];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_B4 = \$techmap2834$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[20].A [3];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_B5 = \counter [12];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_B6 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_BX = \$auto$alumacc.cc:485:replace_alu$1415.Y [12];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_C1 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_C2 = \counter [13];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_C3 = \$techmap2843$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[13].A [2];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_C4 = \counter [12];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_C5 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_C6 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_CX = \$auto$alumacc.cc:485:replace_alu$1415.Y [16];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_D1 = CLBLL_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLL_R_X17Y130_SLICE_X26Y130_D2 = \counter [14];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_D3 = \$techmap2812$abc$2783$lut$aiger2782$119.A [2];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_D4 = \counter [15];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_D5 = \$techmap2812$abc$2783$lut$aiger2782$119.A [3];
  assign CLBLL_R_X17Y130_SLICE_X26Y130_D6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_D3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A2 = CLBLL_R_X17Y120_SLICE_X27Y120_CQ;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A4 = CLBLL_R_X17Y130_SLICE_X27Y130_BO6;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A5 = CLBLL_R_X17Y120_SLICE_X27Y120_C5Q;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_D4 = \$techmap2812$abc$2783$lut$aiger2782$119.A [2];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_D5 = \$techmap2812$abc$2783$lut$aiger2782$119.A [3];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B1 = CLBLL_R_X17Y120_SLICE_X27Y120_CQ;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B2 = CLBLL_R_X17Y120_SLICE_X27Y120_DQ;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B3 = CLBLL_R_X17Y120_SLICE_X27Y120_D5Q;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B4 = CLBLL_R_X17Y130_SLICE_X27Y130_BO6;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B5 = CLBLL_R_X17Y120_SLICE_X27Y120_C5Q;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_D6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C1 = \$auto$alumacc.cc:485:replace_alu$1415.Y [32];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C2 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_A1 = \counter [22];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_A2 = \$techmap2810$abc$2783$lut$aiger2782$176.A [4];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_A3 = \counter [23];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_A4 = \counter [21];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_CX = \$auto$alumacc.cc:485:replace_alu$1415.Y [33];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_A5 = \counter [20];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D2 = \$auto$alumacc.cc:485:replace_alu$1415.Y [34];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D6 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_A6 = \$techmap2810$abc$2783$lut$aiger2782$176.A [5];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_DX = \$auto$alumacc.cc:485:replace_alu$1415.Y [35];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_B1 = \counter [25];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_B2 = CLBLL_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_B3 = \$techmap2813$abc$2783$lut$aiger2782$231.A [2];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_B4 = CLBLL_R_X17Y130_SLICE_X27Y130_AO6;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_B5 = \counter [24];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_B6 = \$techmap2813$abc$2783$lut$aiger2782$231.A [5];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_C1 = \counter [19];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_C2 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_C3 = \$techmap2834$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[20].A [3];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_C4 = \counter [18];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_C5 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_C6 = 1'b1;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_D = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_D = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_CX = \$auto$alumacc.cc:485:replace_alu$1415.Y [18];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_D1 = \counter [21];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_D2 = \counter [20];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_D3 = \$techmap2810$abc$2783$lut$aiger2782$176.A [5];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_D4 = \$techmap2810$abc$2783$lut$aiger2782$176.A [4];
  assign CLBLL_R_X17Y130_SLICE_X27Y130_D5 = CLBLL_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLL_R_X17Y130_SLICE_X27Y130_D6 = \$techmap2813$abc$2783$lut$aiger2782$231.A [5];
  assign RIOI3_X43Y61_OLOGIC_X1Y61_D1 = CLBLL_R_X17Y128_SLICE_X26Y128_BQ;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_T1 = 1'b1;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_D1 = CLBLL_R_X17Y129_SLICE_X26Y129_C5Q;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_T1 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_D1 = CLBLL_R_X17Y120_SLICE_X27Y120_D5Q;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_D1 = CLBLL_R_X17Y120_SLICE_X27Y120_C5Q;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_T1 = 1'b1;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_T1 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_D1 = CLBLL_R_X17Y120_SLICE_X27Y120_DQ;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_T1 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X18Y135_A1 = \counter [7];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_A2 = \counter [6];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_A3 = \counter [3];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_A4 = \counter [4];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_A5 = \counter [5];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_A6 = \$techmap2792$abc$2783$lut$aiger2782$78.A [5];
  assign RIOB33_X43Y61_IOB_X1Y61_O = CLBLL_R_X17Y128_SLICE_X26Y128_BQ;
  assign CLBLL_R_X13Y135_SLICE_X18Y135_B1 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X18Y135_B2 = \counter [1];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_B3 = \counter [7];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_B4 = \$techmap2798$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[6].A [1];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_B5 = \counter [0];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_B6 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X18Y135_BX = \$auto$alumacc.cc:485:replace_alu$1415.Y [5];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_C1 = \counter [2];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_C2 = \counter [0];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_C3 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X18Y135_C4 = \counter [1];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_C5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [7];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_C6 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X18Y135_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X13Y135_SLICE_X18Y135_CX = \$auto$alumacc.cc:485:replace_alu$1415.Y [3];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_D1 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X18Y135_D2 = \counter [3];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_D3 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X18Y135_D4 = \$techmap2792$abc$2783$lut$aiger2782$78.A [5];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_D5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [2];
  assign CLBLL_R_X13Y135_SLICE_X18Y135_D6 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X18Y135_DX = \$auto$alumacc.cc:485:replace_alu$1415.Y [6];
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_D1 = CLBLL_R_X17Y128_SLICE_X26Y128_DQ;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_A1 = \counter [12];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_A2 = \counter [14];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_A3 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_A4 = \$techmap2812$abc$2783$lut$aiger2782$119.A [2];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_A5 = \$techmap2843$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[13].A [2];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_A6 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X19Y135_A1 = \$techmap2797$abc$2783$lut$aiger2782$68.A [3];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_A2 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X19Y135_A3 = \counter [4];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_A4 = \counter [5];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_A5 = \counter [6];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_A6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_B1 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_B2 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_B3 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X19Y135_B1 = \$techmap2797$abc$2783$lut$aiger2782$68.A [3];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_B2 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X19Y135_B3 = \counter [5];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_B4 = \counter [6];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_B5 = \counter [4];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_B6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_B4 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_B5 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X19Y135_C1 = \$techmap2792$abc$2783$lut$aiger2782$78.A [5];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_C2 = \counter [3];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_C3 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X19Y135_C4 = \$auto$alumacc.cc:485:replace_alu$1415.Y [4];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_C5 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X19Y135_C6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_C4 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_C5 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X19Y135_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_D1 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_D2 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_D3 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X19Y135_CX = \$auto$alumacc.cc:485:replace_alu$1415.X [0];
  assign CLBLL_R_X17Y131_SLICE_X26Y131_D4 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X19Y135_D1 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X19Y135_D2 = 1'b1;
  assign CLBLL_R_X13Y135_SLICE_X19Y135_D3 = \counter [0];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_D4 = \counter [2];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_D5 = \counter [1];
  assign CLBLL_R_X13Y135_SLICE_X19Y135_D6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_D5 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X26Y131_D6 = 1'b1;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_D = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_A1 = \$techmap2829$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[23].A [1];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_A2 = \counter [23];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_A3 = \counter [22];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_A4 = CLBLL_R_X17Y130_SLICE_X27Y130_DO6;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_A5 = \counter [24];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_A6 = 1'b1;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_D = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_B1 = \counter [22];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_B2 = CLBLL_R_X17Y130_SLICE_X27Y130_DO6;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_B3 = CLBLL_R_X17Y130_SLICE_X27Y130_AO6;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_B4 = \$techmap2813$abc$2783$lut$aiger2782$231.A [5];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_B5 = CLBLL_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_B6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_C1 = \$techmap2813$abc$2783$lut$aiger2782$231.A [5];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_C2 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_C3 = CLBLL_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_C4 = \$auto$alumacc.cc:485:replace_alu$1415.Y [23];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_A1 = CLBLL_R_X17Y128_SLICE_X26Y128_C5Q;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_A2 = CLBLL_R_X17Y128_SLICE_X26Y128_DQ;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_A3 = CLBLL_R_X17Y128_SLICE_X26Y128_BQ;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_A4 = \counter [25];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_A5 = \$techmap2807$abc$2783$lut$aiger2782$226.A [2];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_A6 = \$techmap2822$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[29].A [5];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_C5 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_C6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_B1 = \$techmap2822$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[29].A [5];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_B2 = \counter [25];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_B3 = \counter [27];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_B4 = \counter [26];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_B5 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_B6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_CX = \$auto$alumacc.cc:485:replace_alu$1415.Y [24];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_D1 = \counter [14];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_BX = \$auto$alumacc.cc:485:replace_alu$1415.Y [28];
  assign CLBLL_R_X17Y131_SLICE_X27Y131_D2 = \counter [15];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_C1 = \$techmap2822$abc$2783$lut$auto$alumacc.cc:485:replace_alu$1415.Y[29].A [5];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_C2 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_C3 = CLBLL_R_X17Y128_SLICE_X26Y128_AO6;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_C4 = \counter [26];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_C5 = \counter [25];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_C6 = 1'b1;
  assign CLBLL_R_X17Y131_SLICE_X27Y131_DX = \$auto$alumacc.cc:485:replace_alu$1415.Y [22];
  assign RIOB33_X43Y55_IOB_X1Y55_O = CLBLL_R_X17Y128_SLICE_X26Y128_C5Q;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_CX = \$auto$alumacc.cc:485:replace_alu$1415.Y [27];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D1 = CLBLL_R_X17Y128_SLICE_X26Y128_BQ;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D2 = CLBLL_R_X17Y128_SLICE_X26Y128_C5Q;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D3 = CLBLL_R_X17Y128_SLICE_X26Y128_DQ;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D4 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [26];
  assign CLBLL_R_X17Y128_SLICE_X26Y128_D6 = 1'b1;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_D1 = CLBLL_R_X17Y120_SLICE_X27Y120_CQ;
  assign CLBLL_R_X17Y128_SLICE_X26Y128_DX = CLBLL_R_X17Y129_SLICE_X27Y129_DO6;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_T1 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_A1 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_A2 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_A3 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_A4 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_A5 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_A6 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_B1 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_B2 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_B3 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_B4 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_B5 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_B6 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_C1 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_C2 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_C3 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_C4 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_C5 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_C6 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_D1 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_D2 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_D3 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_D4 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_D5 = 1'b1;
  assign CLBLL_R_X17Y128_SLICE_X27Y128_D6 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I0 = RIOB33_X43Y75_IOB_X1Y76_I;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I1 = 1'b1;
  assign CLBLL_R_X17Y132_SLICE_X27Y132_D3 = \counter [11];
endmodule
