module top(
  input clk,
  input [7:0] sw,
  output [7:0] led
  );
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A1;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A2;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A3;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A4;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_AO5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_AO6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A_CY;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A_XOR;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B1;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B2;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B3;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B4;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_BO5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_BO6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B_CY;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B_XOR;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C1;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C2;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C3;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C4;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_CO5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_CO6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C_CY;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C_XOR;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D1;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D2;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D3;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D4;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_DO5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_DO6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D_CY;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D_XOR;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A1;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A2;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A3;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A4;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_AMUX;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_AO5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_AO6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_AQ;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_AX;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A_CY;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A_XOR;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B1;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B2;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B3;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B4;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_BMUX;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_BO5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_BO6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_BQ;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_BX;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B_CY;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B_XOR;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C1;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C2;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C3;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C4;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_CLK;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_CMUX;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_CO5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_CO6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_COUT;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_CQ;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_CX;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C_CY;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C_XOR;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D1;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D2;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D3;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D4;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_DMUX;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_DO5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_DO6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_DQ;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_DX;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D_CY;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D_XOR;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A1;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A2;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A3;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A4;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_AO5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_AO6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A_CY;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A_XOR;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B1;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B2;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B3;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B4;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_BO5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_BO6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B_CY;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B_XOR;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C1;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C2;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C3;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C4;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_CO5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_CO6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C_CY;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C_XOR;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D1;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D2;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D3;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D4;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_DO5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_DO6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D_CY;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D_XOR;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A1;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A2;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A3;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A4;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_AMUX;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_AO5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_AO6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_AQ;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_AX;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A_CY;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A_XOR;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B1;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B2;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B3;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B4;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_BMUX;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_BO5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_BO6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_BQ;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_BX;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B_CY;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B_XOR;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C1;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C2;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C3;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C4;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_CIN;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_CLK;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_CMUX;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_CO5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_CO6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_COUT;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_CQ;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_CX;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C_CY;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C_XOR;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D1;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D2;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D3;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D4;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_DMUX;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_DO5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_DO6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_DQ;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_DX;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D_CY;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_AO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_AO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_BO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_BO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_CO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_CO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_DO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_DO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_AO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_AO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_AQ;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_AX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_BMUX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_BO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_BO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_BQ;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_BX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CIN;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CLK;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CMUX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_COUT;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CQ;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_DMUX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_DO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_DO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_DQ;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_DX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D_XOR;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A1;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A2;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A3;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A4;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_AO5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_AO6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A_CY;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A_XOR;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B1;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B2;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B3;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B4;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_BO5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_BO6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B_CY;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B_XOR;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C1;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C2;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C3;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C4;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_CO5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_CO6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C_CY;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C_XOR;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D1;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D2;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D3;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D4;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_DO5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_DO6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D_CY;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D_XOR;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A1;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A2;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A3;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A4;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_AO5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_AO6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_AQ;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_AX;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A_CY;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A_XOR;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B1;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B2;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B3;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B4;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_BMUX;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_BO5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_BO6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_BQ;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_BX;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B_CY;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B_XOR;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C1;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C2;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C3;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C4;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_CIN;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_CLK;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_CMUX;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_CO5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_CO6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_COUT;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_CQ;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_CX;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C_CY;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C_XOR;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D1;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D2;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D3;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D4;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_DMUX;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_DO5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_DO6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_DQ;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_DX;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D_CY;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D_XOR;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S1;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_CE;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_I;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_I;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_O;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y2_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_TQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_TQ;
  wire [0:0] RIOB33_SING_X43Y50_IOB_X1Y50_O;
  wire [0:0] RIOB33_X43Y51_IOB_X1Y51_O;
  wire [0:0] RIOB33_X43Y51_IOB_X1Y52_O;
  wire [0:0] RIOB33_X43Y55_IOB_X1Y55_O;
  wire [0:0] RIOB33_X43Y57_IOB_X1Y58_O;
  wire [0:0] RIOB33_X43Y61_IOB_X1Y61_O;
  wire [0:0] RIOB33_X43Y75_IOB_X1Y76_I;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_D1;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_OQ;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_T1;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_TQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_D1;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_OQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_T1;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_TQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_D1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_OQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_T1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_TQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_D1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_OQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_T1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_TQ;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_D1;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_OQ;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_T1;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_TQ;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_D1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_OQ;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_T1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_TQ;
  wire [0:0] RIOI3_X43Y75_ILOGIC_X1Y76_D;
  wire [0:0] RIOI3_X43Y75_ILOGIC_X1Y76_O;
  wire [0:0] \$abc$3464$aiger3463$35 ;
  wire [0:0] \$abc$3464$aiger3463$44 ;
  wire [0:0] \$abc$3464$aiger3463$53 ;
  wire [15:0] \$auto$alumacc.cc:485:replace_alu$1385.O ;
  wire [7:0] \counter ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y118_SLICE_X26Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y118_SLICE_X26Y118_DO5),
.O6(CLBLL_R_X17Y118_SLICE_X26Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y118_SLICE_X26Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y118_SLICE_X26Y118_CO5),
.O6(CLBLL_R_X17Y118_SLICE_X26Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y118_SLICE_X26Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y118_SLICE_X26Y118_BO5),
.O6(CLBLL_R_X17Y118_SLICE_X26Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y118_SLICE_X26Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y118_SLICE_X26Y118_AO5),
.O6(CLBLL_R_X17Y118_SLICE_X26Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1473CLBLL_R_X17Y118_SLICE_X27Y118_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y118_SLICE_X27Y118_AO5),
.Q(\counter [2]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1474CLBLL_R_X17Y118_SLICE_X27Y118_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y118_SLICE_X27Y118_BO5),
.Q(\counter [3]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1472CLBLL_R_X17Y118_SLICE_X27Y118_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y118_SLICE_X27Y118_CO5),
.Q(\counter [1]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1471CLBLL_R_X17Y118_SLICE_X27Y118_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y118_SLICE_X27Y118_DO5),
.Q(\counter [0]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y118_SLICE_X27Y118_CARRY4 (
.CI(1'b0),
.CO({\$abc$3464$aiger3463$35 , CLBLL_R_X17Y118_SLICE_X27Y118_C_CY, CLBLL_R_X17Y118_SLICE_X27Y118_B_CY, CLBLL_R_X17Y118_SLICE_X27Y118_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({\$auto$alumacc.cc:485:replace_alu$1385.O [3], \$auto$alumacc.cc:485:replace_alu$1385.O [2], \$auto$alumacc.cc:485:replace_alu$1385.O [1], CLBLL_R_X17Y118_SLICE_X27Y118_A_XOR}),
.S({CLBLL_R_X17Y118_SLICE_X27Y118_DO6, CLBLL_R_X17Y118_SLICE_X27Y118_CO6, CLBLL_R_X17Y118_SLICE_X27Y118_BO6, CLBLL_R_X17Y118_SLICE_X27Y118_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLL_R_X17Y118_SLICE_X27Y118_DLUT (
.I0(CLBLL_R_X17Y118_SLICE_X27Y118_AO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(\counter [3]),
.I5(1'b1),
.O5(CLBLL_R_X17Y118_SLICE_X27Y118_DO5),
.O6(CLBLL_R_X17Y118_SLICE_X27Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacccccccc)
  ) CLBLL_R_X17Y118_SLICE_X27Y118_CLUT (
.I0(\counter [2]),
.I1(\$auto$alumacc.cc:485:replace_alu$1385.O [1]),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y118_SLICE_X27Y118_CO5),
.O6(CLBLL_R_X17Y118_SLICE_X27Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y118_SLICE_X27Y118_BLUT (
.I0(1'b1),
.I1(\counter [1]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1385.O [3]),
.I5(1'b1),
.O5(CLBLL_R_X17Y118_SLICE_X27Y118_BO5),
.O6(CLBLL_R_X17Y118_SLICE_X27Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffffff0000)
  ) CLBLL_R_X17Y118_SLICE_X27Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(\counter [0]),
.I4(\$auto$alumacc.cc:485:replace_alu$1385.O [2]),
.I5(1'b1),
.O5(CLBLL_R_X17Y118_SLICE_X27Y118_AO5),
.O6(CLBLL_R_X17Y118_SLICE_X27Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y119_SLICE_X26Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y119_SLICE_X26Y119_DO5),
.O6(CLBLL_R_X17Y119_SLICE_X26Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y119_SLICE_X26Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y119_SLICE_X26Y119_CO5),
.O6(CLBLL_R_X17Y119_SLICE_X26Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y119_SLICE_X26Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y119_SLICE_X26Y119_BO5),
.O6(CLBLL_R_X17Y119_SLICE_X26Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y119_SLICE_X26Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y119_SLICE_X26Y119_AO5),
.O6(CLBLL_R_X17Y119_SLICE_X26Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1477CLBLL_R_X17Y119_SLICE_X27Y119_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y119_SLICE_X27Y119_AO5),
.Q(\counter [6]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1478CLBLL_R_X17Y119_SLICE_X27Y119_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y119_SLICE_X27Y119_BO5),
.Q(\counter [7]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1475CLBLL_R_X17Y119_SLICE_X27Y119_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y119_SLICE_X27Y119_CO5),
.Q(\counter [4]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1476CLBLL_R_X17Y119_SLICE_X27Y119_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y119_SLICE_X27Y119_DO5),
.Q(\counter [5]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y119_SLICE_X27Y119_CARRY4 (
.CI(\$abc$3464$aiger3463$35 ),
.CO({\$abc$3464$aiger3463$44 , CLBLL_R_X17Y119_SLICE_X27Y119_C_CY, CLBLL_R_X17Y119_SLICE_X27Y119_B_CY, CLBLL_R_X17Y119_SLICE_X27Y119_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1385.O [7], \$auto$alumacc.cc:485:replace_alu$1385.O [6], \$auto$alumacc.cc:485:replace_alu$1385.O [5], \$auto$alumacc.cc:485:replace_alu$1385.O [4]}),
.S({CLBLL_R_X17Y119_SLICE_X27Y119_DO6, CLBLL_R_X17Y119_SLICE_X27Y119_CO6, CLBLL_R_X17Y119_SLICE_X27Y119_BO6, CLBLL_R_X17Y119_SLICE_X27Y119_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLL_R_X17Y119_SLICE_X27Y119_DLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1385.O [5]),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(\counter [7]),
.I5(1'b1),
.O5(CLBLL_R_X17Y119_SLICE_X27Y119_DO5),
.O6(CLBLL_R_X17Y119_SLICE_X27Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_R_X17Y119_SLICE_X27Y119_CLUT (
.I0(1'b1),
.I1(\$auto$alumacc.cc:485:replace_alu$1385.O [4]),
.I2(\counter [6]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y119_SLICE_X27Y119_CO5),
.O6(CLBLL_R_X17Y119_SLICE_X27Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y119_SLICE_X27Y119_BLUT (
.I0(1'b1),
.I1(\counter [5]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1385.O [7]),
.I5(1'b1),
.O5(CLBLL_R_X17Y119_SLICE_X27Y119_BO5),
.O6(CLBLL_R_X17Y119_SLICE_X27Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y119_SLICE_X27Y119_ALUT (
.I0(1'b1),
.I1(\counter [4]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1385.O [6]),
.I5(1'b1),
.O5(CLBLL_R_X17Y119_SLICE_X27Y119_AO5),
.O6(CLBLL_R_X17Y119_SLICE_X27Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y120_SLICE_X26Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X26Y120_DO5),
.O6(CLBLL_R_X17Y120_SLICE_X26Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y120_SLICE_X26Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X26Y120_CO5),
.O6(CLBLL_R_X17Y120_SLICE_X26Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y120_SLICE_X26Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X26Y120_BO5),
.O6(CLBLL_R_X17Y120_SLICE_X26Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y120_SLICE_X26Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X26Y120_AO5),
.O6(CLBLL_R_X17Y120_SLICE_X26Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_A_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y120_SLICE_X27Y120_A_XOR),
.Q(CLBLL_R_X17Y120_SLICE_X27Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_B_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y120_SLICE_X27Y120_BO5),
.Q(CLBLL_R_X17Y120_SLICE_X27Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_C_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y120_SLICE_X27Y120_CO5),
.Q(CLBLL_R_X17Y120_SLICE_X27Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_D_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y120_SLICE_X27Y120_DO5),
.Q(CLBLL_R_X17Y120_SLICE_X27Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y120_SLICE_X27Y120_CARRY4 (
.CI(\$abc$3464$aiger3463$44 ),
.CO({\$abc$3464$aiger3463$53 , CLBLL_R_X17Y120_SLICE_X27Y120_C_CY, CLBLL_R_X17Y120_SLICE_X27Y120_B_CY, CLBLL_R_X17Y120_SLICE_X27Y120_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1385.O [11], \$auto$alumacc.cc:485:replace_alu$1385.O [10], \$auto$alumacc.cc:485:replace_alu$1385.O [9], CLBLL_R_X17Y120_SLICE_X27Y120_A_XOR}),
.S({CLBLL_R_X17Y120_SLICE_X27Y120_DO6, CLBLL_R_X17Y120_SLICE_X27Y120_CO6, CLBLL_R_X17Y120_SLICE_X27Y120_BO6, CLBLL_R_X17Y120_SLICE_X27Y120_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ff00)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_R_X17Y120_SLICE_X27Y120_CQ),
.I3(\$auto$alumacc.cc:485:replace_alu$1385.O [9]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X27Y120_DO5),
.O6(CLBLL_R_X17Y120_SLICE_X27Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_CLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1385.O [11]),
.I1(CLBLL_R_X17Y120_SLICE_X27Y120_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X27Y120_CO5),
.O6(CLBLL_R_X17Y120_SLICE_X27Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X17Y120_SLICE_X27Y120_DQ),
.I2(1'b1),
.I3(\$auto$alumacc.cc:485:replace_alu$1385.O [10]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X27Y120_BO5),
.O6(CLBLL_R_X17Y120_SLICE_X27Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X17Y120_SLICE_X27Y120_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X27Y120_AO5),
.O6(CLBLL_R_X17Y120_SLICE_X27Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y121_SLICE_X26Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y121_SLICE_X26Y121_DO5),
.O6(CLBLL_R_X17Y121_SLICE_X26Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y121_SLICE_X26Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y121_SLICE_X26Y121_CO5),
.O6(CLBLL_R_X17Y121_SLICE_X26Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y121_SLICE_X26Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y121_SLICE_X26Y121_BO5),
.O6(CLBLL_R_X17Y121_SLICE_X26Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y121_SLICE_X26Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y121_SLICE_X26Y121_AO5),
.O6(CLBLL_R_X17Y121_SLICE_X26Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y121_SLICE_X27Y121_A_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y121_SLICE_X27Y121_A_XOR),
.Q(CLBLL_R_X17Y121_SLICE_X27Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y121_SLICE_X27Y121_B_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y121_SLICE_X27Y121_BO5),
.Q(CLBLL_R_X17Y121_SLICE_X27Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y121_SLICE_X27Y121_C_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y121_SLICE_X27Y121_CO5),
.Q(CLBLL_R_X17Y121_SLICE_X27Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y121_SLICE_X27Y121_D_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y121_SLICE_X27Y121_DO5),
.Q(CLBLL_R_X17Y121_SLICE_X27Y121_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y121_SLICE_X27Y121_CARRY4 (
.CI(\$abc$3464$aiger3463$53 ),
.CO({CLBLL_R_X17Y121_SLICE_X27Y121_D_CY, CLBLL_R_X17Y121_SLICE_X27Y121_C_CY, CLBLL_R_X17Y121_SLICE_X27Y121_B_CY, CLBLL_R_X17Y121_SLICE_X27Y121_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1385.O [15], \$auto$alumacc.cc:485:replace_alu$1385.O [14], \$auto$alumacc.cc:485:replace_alu$1385.O [13], CLBLL_R_X17Y121_SLICE_X27Y121_A_XOR}),
.S({CLBLL_R_X17Y121_SLICE_X27Y121_DO6, CLBLL_R_X17Y121_SLICE_X27Y121_CO6, CLBLL_R_X17Y121_SLICE_X27Y121_BO6, CLBLL_R_X17Y121_SLICE_X27Y121_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ff00)
  ) CLBLL_R_X17Y121_SLICE_X27Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_R_X17Y121_SLICE_X27Y121_CQ),
.I3(\$auto$alumacc.cc:485:replace_alu$1385.O [13]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y121_SLICE_X27Y121_DO5),
.O6(CLBLL_R_X17Y121_SLICE_X27Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLL_R_X17Y121_SLICE_X27Y121_CLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1385.O [15]),
.I1(CLBLL_R_X17Y121_SLICE_X27Y121_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y121_SLICE_X27Y121_CO5),
.O6(CLBLL_R_X17Y121_SLICE_X27Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLL_R_X17Y121_SLICE_X27Y121_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X17Y121_SLICE_X27Y121_DQ),
.I2(1'b1),
.I3(\$auto$alumacc.cc:485:replace_alu$1385.O [14]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y121_SLICE_X27Y121_BO5),
.O6(CLBLL_R_X17Y121_SLICE_X27Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLL_R_X17Y121_SLICE_X27Y121_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X17Y121_SLICE_X27Y121_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y121_SLICE_X27Y121_AO5),
.O6(CLBLL_R_X17Y121_SLICE_X27Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X43Y75_IOB_X1Y76_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O),
.O(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y1_OBUF (
.I(CLBLL_R_X17Y121_SLICE_X27Y121_CQ),
.O(led[7])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y2_OBUF (
.I(CLBLL_R_X17Y121_SLICE_X27Y121_BQ),
.O(led[6])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y121_IOB_X0Y122_IBUF (
.I(sw[3]),
.O(LIOB33_X0Y121_IOB_X0Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y123_IOB_X0Y123_IBUF (
.I(sw[2]),
.O(LIOB33_X0Y123_IOB_X0Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y123_IOB_X0Y124_IBUF (
.I(sw[1]),
.O(LIOB33_X0Y123_IOB_X0Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y125_IOB_X0Y125_IBUF (
.I(sw[0]),
.O(LIOB33_X0Y125_IOB_X0Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y125_IOB_X0Y126_IBUF (
.I(sw[7]),
.O(LIOB33_X0Y125_IOB_X0Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y127_IOB_X0Y127_IBUF (
.I(sw[6]),
.O(LIOB33_X0Y127_IOB_X0Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(sw[5]),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y137_IOB_X0Y137_IBUF (
.I(sw[4]),
.O(LIOB33_X0Y137_IOB_X0Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y51_IOB_X1Y51_OBUF (
.I(CLBLL_R_X17Y121_SLICE_X27Y121_AQ),
.O(led[4])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y51_IOB_X1Y52_OBUF (
.I(CLBLL_R_X17Y120_SLICE_X27Y120_CQ),
.O(led[3])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y55_IOB_X1Y55_OBUF (
.I(CLBLL_R_X17Y120_SLICE_X27Y120_BQ),
.O(led[2])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y57_IOB_X1Y58_OBUF (
.I(CLBLL_R_X17Y120_SLICE_X27Y120_DQ),
.O(led[1])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y61_IOB_X1Y61_OBUF (
.I(CLBLL_R_X17Y120_SLICE_X27Y120_AQ),
.O(led[0])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y75_IOB_X1Y76_IBUF (
.I(clk),
.O(RIOB33_X43Y75_IOB_X1Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_SING_X43Y50_IOB_X1Y50_OBUF (
.I(CLBLL_R_X17Y121_SLICE_X27Y121_DQ),
.O(led[5])
  );
  assign CLBLL_R_X17Y118_SLICE_X27Y118_COUT = \$abc$3464$aiger3463$35 ;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_AQ = \counter [2];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_BQ = \counter [3];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_CQ = \counter [1];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_DQ = \counter [0];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_BMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [1];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_CMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [2];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_DMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [3];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_COUT = \$abc$3464$aiger3463$44 ;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_AQ = \counter [6];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_BQ = \counter [7];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_CQ = \counter [4];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_DQ = \counter [5];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_AMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [4];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_BMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [5];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_CMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [6];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_DMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [7];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_COUT = \$abc$3464$aiger3463$53 ;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_BMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [9];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_CMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [10];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_DMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [11];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_BMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [13];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_CMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [14];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_DMUX = \$auto$alumacc.cc:485:replace_alu$1385.O [15];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_B_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [1];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_C_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [2];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [3];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D_CY = \$abc$3464$aiger3463$35 ;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_A_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [4];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_B_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [5];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_C_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [6];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [7];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D_CY = \$abc$3464$aiger3463$44 ;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [9];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [10];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [11];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D_CY = \$abc$3464$aiger3463$53 ;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_B_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [13];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_C_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [14];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D_XOR = \$auto$alumacc.cc:485:replace_alu$1385.O [15];
  assign CLBLL_R_X17Y118_SLICE_X26Y118_A = CLBLL_R_X17Y118_SLICE_X26Y118_AO6;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_B = CLBLL_R_X17Y118_SLICE_X26Y118_BO6;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_C = CLBLL_R_X17Y118_SLICE_X26Y118_CO6;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_D = CLBLL_R_X17Y118_SLICE_X26Y118_DO6;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_A = CLBLL_R_X17Y118_SLICE_X27Y118_AO6;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_B = CLBLL_R_X17Y118_SLICE_X27Y118_BO6;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_C = CLBLL_R_X17Y118_SLICE_X27Y118_CO6;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D = CLBLL_R_X17Y118_SLICE_X27Y118_DO6;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_AMUX = CLBLL_R_X17Y118_SLICE_X27Y118_AO6;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_A = CLBLL_R_X17Y119_SLICE_X26Y119_AO6;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_B = CLBLL_R_X17Y119_SLICE_X26Y119_BO6;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_C = CLBLL_R_X17Y119_SLICE_X26Y119_CO6;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_D = CLBLL_R_X17Y119_SLICE_X26Y119_DO6;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_A = CLBLL_R_X17Y119_SLICE_X27Y119_AO6;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_B = CLBLL_R_X17Y119_SLICE_X27Y119_BO6;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_C = CLBLL_R_X17Y119_SLICE_X27Y119_CO6;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D = CLBLL_R_X17Y119_SLICE_X27Y119_DO6;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A = CLBLL_R_X17Y120_SLICE_X26Y120_AO6;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B = CLBLL_R_X17Y120_SLICE_X26Y120_BO6;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C = CLBLL_R_X17Y120_SLICE_X26Y120_CO6;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D = CLBLL_R_X17Y120_SLICE_X26Y120_DO6;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A = CLBLL_R_X17Y120_SLICE_X27Y120_AO6;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B = CLBLL_R_X17Y120_SLICE_X27Y120_BO6;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C = CLBLL_R_X17Y120_SLICE_X27Y120_CO6;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D = CLBLL_R_X17Y120_SLICE_X27Y120_DO6;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_A = CLBLL_R_X17Y121_SLICE_X26Y121_AO6;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_B = CLBLL_R_X17Y121_SLICE_X26Y121_BO6;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_C = CLBLL_R_X17Y121_SLICE_X26Y121_CO6;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_D = CLBLL_R_X17Y121_SLICE_X26Y121_DO6;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_A = CLBLL_R_X17Y121_SLICE_X27Y121_AO6;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_B = CLBLL_R_X17Y121_SLICE_X27Y121_BO6;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_C = CLBLL_R_X17Y121_SLICE_X27Y121_CO6;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D = CLBLL_R_X17Y121_SLICE_X27Y121_DO6;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_OQ = CLBLL_R_X17Y121_SLICE_X27Y121_BQ;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_TQ = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_OQ = CLBLL_R_X17Y121_SLICE_X27Y121_CQ;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_TQ = 1'b1;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_O = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_O = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_O = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_O = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_OQ = CLBLL_R_X17Y120_SLICE_X27Y120_CQ;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_TQ = 1'b1;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_OQ = CLBLL_R_X17Y121_SLICE_X27Y121_AQ;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_TQ = 1'b1;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_OQ = CLBLL_R_X17Y120_SLICE_X27Y120_BQ;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_TQ = 1'b1;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_OQ = CLBLL_R_X17Y120_SLICE_X27Y120_AQ;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_TQ = 1'b1;
  assign RIOI3_X43Y75_ILOGIC_X1Y76_O = RIOB33_X43Y75_IOB_X1Y76_I;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_OQ = CLBLL_R_X17Y121_SLICE_X27Y121_DQ;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_OQ = CLBLL_R_X17Y120_SLICE_X27Y120_DQ;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_TQ = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C2 = CLBLL_R_X17Y120_SLICE_X27Y120_BQ;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_CIN = \$abc$3464$aiger3463$44 ;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_CE = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_CX = 1'b0;
  assign LIOB33_X0Y1_IOB_X0Y1_O = CLBLL_R_X17Y121_SLICE_X27Y121_CQ;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D2 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D3 = CLBLL_R_X17Y120_SLICE_X27Y120_CQ;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D4 = \$auto$alumacc.cc:485:replace_alu$1385.O [9];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D6 = 1'b1;
  assign LIOB33_X0Y1_IOB_X0Y2_O = CLBLL_R_X17Y121_SLICE_X27Y121_BQ;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_D = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_DX = 1'b0;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_D = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_D = LIOB33_X0Y125_IOB_X0Y125_I;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_D1 = CLBLL_R_X17Y120_SLICE_X27Y120_AQ;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_T1 = 1'b1;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_D = LIOB33_X0Y121_IOB_X0Y122_I;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_D1 = CLBLL_R_X17Y120_SLICE_X27Y120_BQ;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_A1 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_A2 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_A3 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_A4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_A5 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_A6 = 1'b1;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_B1 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_B2 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_B3 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_B4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_B5 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_B6 = 1'b1;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_D1 = CLBLL_R_X17Y120_SLICE_X27Y120_CQ;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_C1 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_C2 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_C3 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_C4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_C5 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_C6 = 1'b1;
  assign RIOB33_X43Y57_IOB_X1Y58_O = CLBLL_R_X17Y120_SLICE_X27Y120_DQ;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_T1 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_D1 = CLBLL_R_X17Y121_SLICE_X27Y121_BQ;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_D1 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_D2 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_D3 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_D4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_D5 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_D6 = 1'b1;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_D1 = CLBLL_R_X17Y121_SLICE_X27Y121_AQ;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_T1 = 1'b1;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_T1 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_D1 = CLBLL_R_X17Y121_SLICE_X27Y121_CQ;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_T1 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_A1 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_A2 = \counter [4];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_A3 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_A4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_A5 = \$auto$alumacc.cc:485:replace_alu$1385.O [6];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_A6 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_AX = 1'b0;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_B1 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_B2 = \counter [5];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_B3 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_B4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_B5 = \$auto$alumacc.cc:485:replace_alu$1385.O [7];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_B6 = 1'b1;
  assign RIOB33_X43Y61_IOB_X1Y61_O = CLBLL_R_X17Y120_SLICE_X27Y120_AQ;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_BX = 1'b0;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_C1 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_C2 = \$auto$alumacc.cc:485:replace_alu$1385.O [4];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_C3 = \counter [6];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_C4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_C5 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_C6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_CIN = \$abc$3464$aiger3463$35 ;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_CX = 1'b0;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D1 = \$auto$alumacc.cc:485:replace_alu$1385.O [5];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D2 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D3 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D5 = \counter [7];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_A1 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_A2 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_DX = 1'b0;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_A3 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_A4 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_A5 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_A6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_B1 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_B2 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_B3 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_B4 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_B5 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_B6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_C1 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_C2 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_C3 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_C4 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_C5 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_D1 = CLBLL_R_X17Y120_SLICE_X27Y120_DQ;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D3 = CLBLL_R_X17Y121_SLICE_X27Y121_CQ;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_T1 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_D1 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_D2 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_D3 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_D4 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_D5 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_D6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D4 = \$auto$alumacc.cc:485:replace_alu$1385.O [13];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D5 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D6 = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_D = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_A1 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_A2 = CLBLL_R_X17Y121_SLICE_X27Y121_AQ;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_A3 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_A4 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_A5 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_A6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_AX = 1'b0;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_B1 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_B2 = CLBLL_R_X17Y121_SLICE_X27Y121_DQ;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_B3 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_B4 = \$auto$alumacc.cc:485:replace_alu$1385.O [14];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_B5 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_B6 = 1'b1;
  assign RIOB33_X43Y51_IOB_X1Y52_O = CLBLL_R_X17Y120_SLICE_X27Y120_CQ;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_BX = 1'b0;
  assign RIOB33_X43Y51_IOB_X1Y51_O = CLBLL_R_X17Y121_SLICE_X27Y121_AQ;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_C1 = \$auto$alumacc.cc:485:replace_alu$1385.O [15];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_C2 = CLBLL_R_X17Y121_SLICE_X27Y121_BQ;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_C3 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_C4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_A1 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_A2 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_A3 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_A4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_A5 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_A6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_C5 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_C6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_CIN = \$abc$3464$aiger3463$53 ;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_B1 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_B2 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_B3 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_B4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_B5 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_B6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_CX = 1'b0;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D1 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D2 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_C1 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_C2 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_C3 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_C4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_C5 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_C6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_DX = 1'b0;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_D1 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_D2 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_D3 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_D4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_D5 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_D6 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE0 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE1 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE0 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE1 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S0 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S1 = 1'b1;
  assign RIOB33_X43Y55_IOB_X1Y55_O = CLBLL_R_X17Y120_SLICE_X27Y120_BQ;
  assign RIOB33_SING_X43Y50_IOB_X1Y50_O = CLBLL_R_X17Y121_SLICE_X27Y121_DQ;
  assign RIOI3_X43Y75_ILOGIC_X1Y76_D = RIOB33_X43Y75_IOB_X1Y76_I;
  assign CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_I = CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_D1 = CLBLL_R_X17Y121_SLICE_X27Y121_DQ;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_A1 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_A2 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_A3 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_A4 = \counter [0];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_A5 = \$auto$alumacc.cc:485:replace_alu$1385.O [2];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_A6 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_AX = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_B1 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_B2 = \counter [1];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_B3 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_B4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_B5 = \$auto$alumacc.cc:485:replace_alu$1385.O [3];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_B6 = 1'b1;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_T1 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_BX = 1'b0;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_C1 = \counter [2];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_C2 = \$auto$alumacc.cc:485:replace_alu$1385.O [1];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_C3 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_C4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_C5 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_C6 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_CX = 1'b0;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D1 = CLBLL_R_X17Y118_SLICE_X27Y118_AO6;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D2 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D3 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D5 = \counter [3];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A2 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_DX = 1'b0;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B2 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C2 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D2 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A2 = CLBLL_R_X17Y120_SLICE_X27Y120_AQ;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_AX = 1'b0;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I0 = RIOB33_X43Y75_IOB_X1Y76_I;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B2 = CLBLL_R_X17Y120_SLICE_X27Y120_DQ;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B4 = \$auto$alumacc.cc:485:replace_alu$1385.O [10];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B6 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I1 = 1'b1;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_D = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_BX = 1'b0;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C1 = \$auto$alumacc.cc:485:replace_alu$1385.O [11];
endmodule
