module top(
  input clk,
  input [7:0] sw,
  output [7:0] led
  );
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_A;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_A1;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_A2;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_A3;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_A4;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_A5;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_A6;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_AO5;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_AO6;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_A_CY;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_A_XOR;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_B;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_B1;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_B2;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_B3;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_B4;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_B5;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_B6;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_BO5;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_BO6;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_B_CY;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_B_XOR;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_C;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_C1;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_C2;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_C3;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_C4;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_C5;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_C6;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_CO5;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_CO6;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_C_CY;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_C_XOR;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_D;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_D1;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_D2;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_D3;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_D4;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_D5;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_D6;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_DO5;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_DO6;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_D_CY;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X26Y115_D_XOR;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_A;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_A1;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_A2;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_A3;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_A4;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_A5;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_A6;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_AO5;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_AO6;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_AQ;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_AX;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_A_CY;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_A_XOR;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_B;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_B1;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_B2;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_B3;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_B4;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_B5;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_B6;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_BMUX;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_BO5;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_BO6;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_BQ;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_BX;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_B_CY;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_B_XOR;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_C;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_C1;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_C2;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_C3;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_C4;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_C5;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_C6;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_CLK;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_CMUX;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_CO5;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_CO6;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_COUT;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_CQ;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_CX;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_C_CY;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_C_XOR;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_D;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_D1;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_D2;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_D3;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_D4;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_D5;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_D6;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_DMUX;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_DO5;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_DO6;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_DQ;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_DX;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_D_CY;
  wire [0:0] CLBLL_R_X17Y115_SLICE_X27Y115_D_XOR;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_A;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_A1;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_A2;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_A3;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_A4;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_A5;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_A6;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_AO5;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_AO6;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_A_CY;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_A_XOR;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_B;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_B1;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_B2;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_B3;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_B4;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_B5;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_B6;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_BO5;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_BO6;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_B_CY;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_B_XOR;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_C;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_C1;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_C2;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_C3;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_C4;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_C5;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_C6;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_CO5;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_CO6;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_C_CY;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_C_XOR;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_D;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_D1;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_D2;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_D3;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_D4;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_D5;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_D6;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_DO5;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_DO6;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_D_CY;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X26Y116_D_XOR;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_A;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_A1;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_A2;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_A3;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_A4;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_A5;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_A6;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_AMUX;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_AO5;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_AO6;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_AQ;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_AX;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_A_CY;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_A_XOR;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_B;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_B1;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_B2;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_B3;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_B4;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_B5;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_B6;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_BMUX;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_BO5;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_BO6;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_BQ;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_BX;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_B_CY;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_B_XOR;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_C;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_C1;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_C2;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_C3;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_C4;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_C5;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_C6;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_CIN;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_CLK;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_CMUX;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_CO5;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_CO6;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_COUT;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_CQ;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_CX;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_C_CY;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_C_XOR;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_D;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_D1;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_D2;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_D3;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_D4;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_D5;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_D6;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_DMUX;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_DO5;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_DO6;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_DQ;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_DX;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_D_CY;
  wire [0:0] CLBLL_R_X17Y116_SLICE_X27Y116_D_XOR;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_A;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_A1;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_A2;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_A3;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_A4;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_A5;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_A6;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_AO5;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_AO6;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_A_CY;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_A_XOR;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_B;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_B1;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_B2;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_B3;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_B4;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_B5;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_B6;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_BO5;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_BO6;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_B_CY;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_B_XOR;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_C;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_C1;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_C2;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_C3;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_C4;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_C5;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_C6;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_CO5;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_CO6;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_C_CY;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_C_XOR;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_D;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_D1;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_D2;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_D3;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_D4;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_D5;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_D6;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_DO5;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_DO6;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_D_CY;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X26Y117_D_XOR;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_A;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_A1;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_A2;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_A3;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_A4;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_A5;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_A6;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_AMUX;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_AO5;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_AO6;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_AQ;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_AX;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_A_CY;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_A_XOR;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_B;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_B1;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_B2;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_B3;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_B4;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_B5;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_B6;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_BMUX;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_BO5;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_BO6;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_BQ;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_BX;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_B_CY;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_B_XOR;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_C;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_C1;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_C2;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_C3;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_C4;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_C5;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_C6;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_CIN;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_CLK;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_CMUX;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_CO5;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_CO6;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_COUT;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_CQ;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_CX;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_C_CY;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_C_XOR;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_D;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_D1;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_D2;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_D3;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_D4;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_D5;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_D6;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_DMUX;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_DO5;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_DO6;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_DQ;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_DX;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_D_CY;
  wire [0:0] CLBLL_R_X17Y117_SLICE_X27Y117_D_XOR;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A1;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A2;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A3;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A4;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_AO5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_AO6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A_CY;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_A_XOR;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B1;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B2;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B3;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B4;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_BO5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_BO6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B_CY;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_B_XOR;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C1;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C2;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C3;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C4;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_CO5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_CO6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C_CY;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_C_XOR;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D1;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D2;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D3;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D4;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_DO5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_DO6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D_CY;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X26Y118_D_XOR;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A1;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A2;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A3;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A4;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_AMUX;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_AO5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_AO6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_AQ;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_AX;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A_CY;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_A_XOR;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B1;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B2;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B3;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B4;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_BMUX;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_BO5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_BO6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_BQ;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_BX;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B_CY;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_B_XOR;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C1;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C2;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C3;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C4;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_CIN;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_CLK;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_CMUX;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_CO5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_CO6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_COUT;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_CQ;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_CX;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C_CY;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_C_XOR;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D1;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D2;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D3;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D4;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_DMUX;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_DO5;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_DO6;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_DQ;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_DX;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D_CY;
  wire [0:0] CLBLL_R_X17Y118_SLICE_X27Y118_D_XOR;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A1;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A2;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A3;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A4;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_AO5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_AO6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A_CY;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_A_XOR;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B1;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B2;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B3;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B4;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_BO5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_BO6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B_CY;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_B_XOR;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C1;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C2;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C3;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C4;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_CO5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_CO6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C_CY;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_C_XOR;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D1;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D2;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D3;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D4;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_DO5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_DO6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D_CY;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X26Y119_D_XOR;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A1;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A2;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A3;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A4;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_AO5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_AO6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_AQ;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_AX;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A_CY;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_A_XOR;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B1;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B2;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B3;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B4;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_BMUX;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_BO5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_BO6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_BQ;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_BX;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B_CY;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_B_XOR;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C1;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C2;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C3;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C4;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_CIN;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_CLK;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_CMUX;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_CO5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_CO6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_COUT;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_CQ;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_CX;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C_CY;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_C_XOR;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D1;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D2;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D3;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D4;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_DMUX;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_DO5;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_DO6;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_DQ;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_DX;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D_CY;
  wire [0:0] CLBLL_R_X17Y119_SLICE_X27Y119_D_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_AO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_AO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_A_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_BO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_BO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_B_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_CO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_CO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_C_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_DO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_DO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X26Y120_D_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_AO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_AO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_AQ;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_AX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_A_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_BMUX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_BO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_BO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_BQ;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_BX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_B_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CIN;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CLK;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CMUX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_COUT;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CQ;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_CX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_C_XOR;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D1;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D2;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D3;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D4;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_DMUX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_DO5;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_DO6;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_DQ;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_DX;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D_CY;
  wire [0:0] CLBLL_R_X17Y120_SLICE_X27Y120_D_XOR;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A1;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A2;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A3;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A4;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_AO5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_AO6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A_CY;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_A_XOR;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B1;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B2;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B3;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B4;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_BO5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_BO6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B_CY;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_B_XOR;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C1;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C2;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C3;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C4;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_CO5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_CO6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C_CY;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_C_XOR;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D1;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D2;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D3;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D4;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_DO5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_DO6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D_CY;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X26Y121_D_XOR;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A1;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A2;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A3;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A4;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_AO5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_AO6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_AQ;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_AX;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A_CY;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_A_XOR;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B1;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B2;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B3;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B4;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_BMUX;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_BO5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_BO6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_BQ;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_BX;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B_CY;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_B_XOR;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C1;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C2;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C3;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C4;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_CIN;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_CLK;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_CMUX;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_CO5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_CO6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_COUT;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_CQ;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_CX;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C_CY;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_C_XOR;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D1;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D2;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D3;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D4;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_DMUX;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_DO5;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_DO6;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_DQ;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_DX;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D_CY;
  wire [0:0] CLBLL_R_X17Y121_SLICE_X27Y121_D_XOR;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_A;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_A1;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_A2;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_A3;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_A4;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_A5;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_A6;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_AO5;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_AO6;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_A_CY;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_A_XOR;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_B;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_B1;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_B2;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_B3;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_B4;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_B5;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_B6;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_BO5;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_BO6;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_B_CY;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_B_XOR;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_C;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_C1;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_C2;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_C3;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_C4;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_C5;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_C6;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_CO5;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_CO6;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_C_CY;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_C_XOR;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_D;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_D1;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_D2;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_D3;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_D4;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_D5;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_D6;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_DO5;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_DO6;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_D_CY;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X26Y122_D_XOR;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_A;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_A1;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_A2;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_A3;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_A4;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_A5;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_A6;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_AO5;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_AO6;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_AQ;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_AX;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_A_CY;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_A_XOR;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_B;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_B1;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_B2;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_B3;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_B4;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_B5;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_B6;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_BMUX;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_BO5;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_BO6;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_BQ;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_BX;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_B_CY;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_B_XOR;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_C;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_C1;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_C2;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_C3;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_C4;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_C5;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_C6;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_CIN;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_CLK;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_CMUX;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_CO5;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_CO6;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_COUT;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_CQ;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_CX;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_C_CY;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_C_XOR;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_D;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_D1;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_D2;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_D3;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_D4;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_D5;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_D6;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_DMUX;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_DO5;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_DO6;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_DQ;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_DX;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_D_CY;
  wire [0:0] CLBLL_R_X17Y122_SLICE_X27Y122_D_XOR;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_A;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_A1;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_A2;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_A3;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_A4;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_A5;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_A6;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_AO5;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_AO6;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_A_CY;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_A_XOR;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_B;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_B1;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_B2;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_B3;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_B4;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_B5;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_B6;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_BO5;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_BO6;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_B_CY;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_B_XOR;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_C;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_C1;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_C2;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_C3;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_C4;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_C5;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_C6;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_CO5;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_CO6;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_C_CY;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_C_XOR;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_D;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_D1;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_D2;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_D3;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_D4;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_D5;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_D6;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_DO5;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_DO6;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_D_CY;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X26Y123_D_XOR;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_A;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_A1;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_A2;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_A3;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_A4;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_A5;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_A6;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_AO5;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_AO6;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_AQ;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_AX;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_A_CY;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_A_XOR;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_B;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_B1;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_B2;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_B3;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_B4;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_B5;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_B6;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_BMUX;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_BO5;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_BO6;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_BQ;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_BX;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_B_CY;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_B_XOR;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_C;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_C1;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_C2;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_C3;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_C4;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_C5;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_C6;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_CIN;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_CLK;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_CMUX;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_CO5;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_CO6;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_COUT;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_CQ;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_CX;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_C_CY;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_C_XOR;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_D;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_D1;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_D2;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_D3;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_D4;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_D5;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_D6;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_DMUX;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_DO5;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_DO6;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_DQ;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_DX;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_D_CY;
  wire [0:0] CLBLL_R_X17Y123_SLICE_X27Y123_D_XOR;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE1;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S0;
  wire [0:0] CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S1;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_CE;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_I;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_I;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_O;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y2_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_TQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_TQ;
  wire [0:0] RIOB33_SING_X43Y50_IOB_X1Y50_O;
  wire [0:0] RIOB33_X43Y51_IOB_X1Y51_O;
  wire [0:0] RIOB33_X43Y51_IOB_X1Y52_O;
  wire [0:0] RIOB33_X43Y55_IOB_X1Y55_O;
  wire [0:0] RIOB33_X43Y57_IOB_X1Y58_O;
  wire [0:0] RIOB33_X43Y61_IOB_X1Y61_O;
  wire [0:0] RIOB33_X43Y75_IOB_X1Y76_I;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_D1;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_OQ;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_T1;
  wire [0:0] RIOI3_SING_X43Y50_OLOGIC_X1Y50_TQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_D1;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_OQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_T1;
  wire [0:0] RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_TQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_D1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_OQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_T1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y51_TQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_D1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_OQ;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_T1;
  wire [0:0] RIOI3_X43Y51_OLOGIC_X1Y52_TQ;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_D1;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_OQ;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_T1;
  wire [0:0] RIOI3_X43Y55_OLOGIC_X1Y55_TQ;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_D1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_OQ;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_T1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_TQ;
  wire [0:0] RIOI3_X43Y75_ILOGIC_X1Y76_D;
  wire [0:0] RIOI3_X43Y75_ILOGIC_X1Y76_O;
  wire [0:0] \$abc$3581$techmap2144$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[1].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  wire [0:0] \$abc$3581$techmap2145$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[2].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  wire [0:0] \$abc$3581$techmap2146$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[3].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  wire [0:0] \$abc$3581$techmap2147$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[4].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  wire [0:0] \$abc$3581$techmap2148$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[5].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  wire [0:0] \$abc$3581$techmap2149$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[6].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  wire [0:0] \$abc$3581$techmap2150$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[7].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  wire [0:0] \$abc$3581$techmap2151$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[8].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  wire [35:0] \$auto$alumacc.cc:485:replace_alu$1415.Y ;
  wire [27:0] \counter ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y115_SLICE_X26Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y115_SLICE_X26Y115_DO5),
.O6(CLBLL_R_X17Y115_SLICE_X26Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y115_SLICE_X26Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y115_SLICE_X26Y115_CO5),
.O6(CLBLL_R_X17Y115_SLICE_X26Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y115_SLICE_X26Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y115_SLICE_X26Y115_BO5),
.O6(CLBLL_R_X17Y115_SLICE_X26Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y115_SLICE_X26Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y115_SLICE_X26Y115_AO5),
.O6(CLBLL_R_X17Y115_SLICE_X26Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1503CLBLL_R_X17Y115_SLICE_X27Y115_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y115_SLICE_X27Y115_AO6),
.Q(\counter [0]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1505CLBLL_R_X17Y115_SLICE_X27Y115_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y115_SLICE_X27Y115_BO5),
.Q(\counter [2]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1506CLBLL_R_X17Y115_SLICE_X27Y115_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y115_SLICE_X27Y115_CO5),
.Q(\counter [3]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1504CLBLL_R_X17Y115_SLICE_X27Y115_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y115_SLICE_X27Y115_DO5),
.Q(\counter [1]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y115_SLICE_X27Y115_CARRY4 (
.CI(1'b0),
.CO({\$abc$3581$techmap2144$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[1].genblk1.carry4.genblk2.genblk1.cin_from_below , CLBLL_R_X17Y115_SLICE_X27Y115_C_CY, CLBLL_R_X17Y115_SLICE_X27Y115_B_CY, CLBLL_R_X17Y115_SLICE_X27Y115_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({\$auto$alumacc.cc:485:replace_alu$1415.Y [3], \$auto$alumacc.cc:485:replace_alu$1415.Y [2], \$auto$alumacc.cc:485:replace_alu$1415.Y [1], CLBLL_R_X17Y115_SLICE_X27Y115_A_XOR}),
.S({CLBLL_R_X17Y115_SLICE_X27Y115_DO6, CLBLL_R_X17Y115_SLICE_X27Y115_CO6, CLBLL_R_X17Y115_SLICE_X27Y115_BO6, CLBLL_R_X17Y115_SLICE_X27Y115_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff00ff00)
  ) CLBLL_R_X17Y115_SLICE_X27Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(\$auto$alumacc.cc:485:replace_alu$1415.Y [1]),
.I4(\counter [3]),
.I5(1'b1),
.O5(CLBLL_R_X17Y115_SLICE_X27Y115_DO5),
.O6(CLBLL_R_X17Y115_SLICE_X27Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaaaaaaa)
  ) CLBLL_R_X17Y115_SLICE_X27Y115_CLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1415.Y [3]),
.I1(1'b1),
.I2(\counter [2]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y115_SLICE_X27Y115_CO5),
.O6(CLBLL_R_X17Y115_SLICE_X27Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0f0f0f0)
  ) CLBLL_R_X17Y115_SLICE_X27Y115_BLUT (
.I0(1'b1),
.I1(\counter [1]),
.I2(\$auto$alumacc.cc:485:replace_alu$1415.Y [2]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y115_SLICE_X27Y115_BO5),
.O6(CLBLL_R_X17Y115_SLICE_X27Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00000000)
  ) CLBLL_R_X17Y115_SLICE_X27Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(\counter [0]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y115_SLICE_X27Y115_AO5),
.O6(CLBLL_R_X17Y115_SLICE_X27Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y116_SLICE_X26Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y116_SLICE_X26Y116_DO5),
.O6(CLBLL_R_X17Y116_SLICE_X26Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y116_SLICE_X26Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y116_SLICE_X26Y116_CO5),
.O6(CLBLL_R_X17Y116_SLICE_X26Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y116_SLICE_X26Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y116_SLICE_X26Y116_BO5),
.O6(CLBLL_R_X17Y116_SLICE_X26Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y116_SLICE_X26Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y116_SLICE_X26Y116_AO5),
.O6(CLBLL_R_X17Y116_SLICE_X26Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1509CLBLL_R_X17Y116_SLICE_X27Y116_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y116_SLICE_X27Y116_AO5),
.Q(\counter [6]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1510CLBLL_R_X17Y116_SLICE_X27Y116_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y116_SLICE_X27Y116_BO5),
.Q(\counter [7]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1507CLBLL_R_X17Y116_SLICE_X27Y116_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y116_SLICE_X27Y116_CO5),
.Q(\counter [4]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1508CLBLL_R_X17Y116_SLICE_X27Y116_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y116_SLICE_X27Y116_DO5),
.Q(\counter [5]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y116_SLICE_X27Y116_CARRY4 (
.CI(\$abc$3581$techmap2144$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[1].genblk1.carry4.genblk2.genblk1.cin_from_below ),
.CO({\$abc$3581$techmap2145$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[2].genblk1.carry4.genblk2.genblk1.cin_from_below , CLBLL_R_X17Y116_SLICE_X27Y116_C_CY, CLBLL_R_X17Y116_SLICE_X27Y116_B_CY, CLBLL_R_X17Y116_SLICE_X27Y116_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1415.Y [7], \$auto$alumacc.cc:485:replace_alu$1415.Y [6], \$auto$alumacc.cc:485:replace_alu$1415.Y [5], \$auto$alumacc.cc:485:replace_alu$1415.Y [4]}),
.S({CLBLL_R_X17Y116_SLICE_X27Y116_DO6, CLBLL_R_X17Y116_SLICE_X27Y116_CO6, CLBLL_R_X17Y116_SLICE_X27Y116_BO6, CLBLL_R_X17Y116_SLICE_X27Y116_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLL_R_X17Y116_SLICE_X27Y116_DLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1415.Y [5]),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(\counter [7]),
.I5(1'b1),
.O5(CLBLL_R_X17Y116_SLICE_X27Y116_DO5),
.O6(CLBLL_R_X17Y116_SLICE_X27Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_R_X17Y116_SLICE_X27Y116_CLUT (
.I0(1'b1),
.I1(\$auto$alumacc.cc:485:replace_alu$1415.Y [4]),
.I2(\counter [6]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y116_SLICE_X27Y116_CO5),
.O6(CLBLL_R_X17Y116_SLICE_X27Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y116_SLICE_X27Y116_BLUT (
.I0(1'b1),
.I1(\counter [5]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1415.Y [7]),
.I5(1'b1),
.O5(CLBLL_R_X17Y116_SLICE_X27Y116_BO5),
.O6(CLBLL_R_X17Y116_SLICE_X27Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y116_SLICE_X27Y116_ALUT (
.I0(1'b1),
.I1(\counter [4]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1415.Y [6]),
.I5(1'b1),
.O5(CLBLL_R_X17Y116_SLICE_X27Y116_AO5),
.O6(CLBLL_R_X17Y116_SLICE_X27Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y117_SLICE_X26Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y117_SLICE_X26Y117_DO5),
.O6(CLBLL_R_X17Y117_SLICE_X26Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y117_SLICE_X26Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y117_SLICE_X26Y117_CO5),
.O6(CLBLL_R_X17Y117_SLICE_X26Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y117_SLICE_X26Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y117_SLICE_X26Y117_BO5),
.O6(CLBLL_R_X17Y117_SLICE_X26Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y117_SLICE_X26Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y117_SLICE_X26Y117_AO5),
.O6(CLBLL_R_X17Y117_SLICE_X26Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1513CLBLL_R_X17Y117_SLICE_X27Y117_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y117_SLICE_X27Y117_AO5),
.Q(\counter [10]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1514CLBLL_R_X17Y117_SLICE_X27Y117_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y117_SLICE_X27Y117_BO5),
.Q(\counter [11]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1511CLBLL_R_X17Y117_SLICE_X27Y117_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y117_SLICE_X27Y117_CO5),
.Q(\counter [8]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1512CLBLL_R_X17Y117_SLICE_X27Y117_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y117_SLICE_X27Y117_DO5),
.Q(\counter [9]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y117_SLICE_X27Y117_CARRY4 (
.CI(\$abc$3581$techmap2145$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[2].genblk1.carry4.genblk2.genblk1.cin_from_below ),
.CO({\$abc$3581$techmap2146$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[3].genblk1.carry4.genblk2.genblk1.cin_from_below , CLBLL_R_X17Y117_SLICE_X27Y117_C_CY, CLBLL_R_X17Y117_SLICE_X27Y117_B_CY, CLBLL_R_X17Y117_SLICE_X27Y117_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1415.Y [11], \$auto$alumacc.cc:485:replace_alu$1415.Y [10], \$auto$alumacc.cc:485:replace_alu$1415.Y [9], \$auto$alumacc.cc:485:replace_alu$1415.Y [8]}),
.S({CLBLL_R_X17Y117_SLICE_X27Y117_DO6, CLBLL_R_X17Y117_SLICE_X27Y117_CO6, CLBLL_R_X17Y117_SLICE_X27Y117_BO6, CLBLL_R_X17Y117_SLICE_X27Y117_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLL_R_X17Y117_SLICE_X27Y117_DLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1415.Y [9]),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(\counter [11]),
.I5(1'b1),
.O5(CLBLL_R_X17Y117_SLICE_X27Y117_DO5),
.O6(CLBLL_R_X17Y117_SLICE_X27Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_R_X17Y117_SLICE_X27Y117_CLUT (
.I0(1'b1),
.I1(\$auto$alumacc.cc:485:replace_alu$1415.Y [8]),
.I2(\counter [10]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y117_SLICE_X27Y117_CO5),
.O6(CLBLL_R_X17Y117_SLICE_X27Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y117_SLICE_X27Y117_BLUT (
.I0(1'b1),
.I1(\counter [9]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1415.Y [11]),
.I5(1'b1),
.O5(CLBLL_R_X17Y117_SLICE_X27Y117_BO5),
.O6(CLBLL_R_X17Y117_SLICE_X27Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y117_SLICE_X27Y117_ALUT (
.I0(1'b1),
.I1(\counter [8]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1415.Y [10]),
.I5(1'b1),
.O5(CLBLL_R_X17Y117_SLICE_X27Y117_AO5),
.O6(CLBLL_R_X17Y117_SLICE_X27Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y118_SLICE_X26Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y118_SLICE_X26Y118_DO5),
.O6(CLBLL_R_X17Y118_SLICE_X26Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y118_SLICE_X26Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y118_SLICE_X26Y118_CO5),
.O6(CLBLL_R_X17Y118_SLICE_X26Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y118_SLICE_X26Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y118_SLICE_X26Y118_BO5),
.O6(CLBLL_R_X17Y118_SLICE_X26Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y118_SLICE_X26Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y118_SLICE_X26Y118_AO5),
.O6(CLBLL_R_X17Y118_SLICE_X26Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1517CLBLL_R_X17Y118_SLICE_X27Y118_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y118_SLICE_X27Y118_AO5),
.Q(\counter [14]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1518CLBLL_R_X17Y118_SLICE_X27Y118_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y118_SLICE_X27Y118_BO5),
.Q(\counter [15]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1515CLBLL_R_X17Y118_SLICE_X27Y118_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y118_SLICE_X27Y118_CO5),
.Q(\counter [12]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1516CLBLL_R_X17Y118_SLICE_X27Y118_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y118_SLICE_X27Y118_DO5),
.Q(\counter [13]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y118_SLICE_X27Y118_CARRY4 (
.CI(\$abc$3581$techmap2146$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[3].genblk1.carry4.genblk2.genblk1.cin_from_below ),
.CO({\$abc$3581$techmap2147$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[4].genblk1.carry4.genblk2.genblk1.cin_from_below , CLBLL_R_X17Y118_SLICE_X27Y118_C_CY, CLBLL_R_X17Y118_SLICE_X27Y118_B_CY, CLBLL_R_X17Y118_SLICE_X27Y118_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1415.Y [15], \$auto$alumacc.cc:485:replace_alu$1415.Y [14], \$auto$alumacc.cc:485:replace_alu$1415.Y [13], \$auto$alumacc.cc:485:replace_alu$1415.Y [12]}),
.S({CLBLL_R_X17Y118_SLICE_X27Y118_DO6, CLBLL_R_X17Y118_SLICE_X27Y118_CO6, CLBLL_R_X17Y118_SLICE_X27Y118_BO6, CLBLL_R_X17Y118_SLICE_X27Y118_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLL_R_X17Y118_SLICE_X27Y118_DLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1415.Y [13]),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(\counter [15]),
.I5(1'b1),
.O5(CLBLL_R_X17Y118_SLICE_X27Y118_DO5),
.O6(CLBLL_R_X17Y118_SLICE_X27Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_R_X17Y118_SLICE_X27Y118_CLUT (
.I0(1'b1),
.I1(\$auto$alumacc.cc:485:replace_alu$1415.Y [12]),
.I2(\counter [14]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y118_SLICE_X27Y118_CO5),
.O6(CLBLL_R_X17Y118_SLICE_X27Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y118_SLICE_X27Y118_BLUT (
.I0(1'b1),
.I1(\counter [13]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1415.Y [15]),
.I5(1'b1),
.O5(CLBLL_R_X17Y118_SLICE_X27Y118_BO5),
.O6(CLBLL_R_X17Y118_SLICE_X27Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y118_SLICE_X27Y118_ALUT (
.I0(1'b1),
.I1(\counter [12]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1415.Y [14]),
.I5(1'b1),
.O5(CLBLL_R_X17Y118_SLICE_X27Y118_AO5),
.O6(CLBLL_R_X17Y118_SLICE_X27Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y119_SLICE_X26Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y119_SLICE_X26Y119_DO5),
.O6(CLBLL_R_X17Y119_SLICE_X26Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y119_SLICE_X26Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y119_SLICE_X26Y119_CO5),
.O6(CLBLL_R_X17Y119_SLICE_X26Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y119_SLICE_X26Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y119_SLICE_X26Y119_BO5),
.O6(CLBLL_R_X17Y119_SLICE_X26Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y119_SLICE_X26Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y119_SLICE_X26Y119_AO5),
.O6(CLBLL_R_X17Y119_SLICE_X26Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1519CLBLL_R_X17Y119_SLICE_X27Y119_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y119_SLICE_X27Y119_A_XOR),
.Q(\counter [16]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1521CLBLL_R_X17Y119_SLICE_X27Y119_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y119_SLICE_X27Y119_BO5),
.Q(\counter [18]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1522CLBLL_R_X17Y119_SLICE_X27Y119_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y119_SLICE_X27Y119_CO5),
.Q(\counter [19]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1520CLBLL_R_X17Y119_SLICE_X27Y119_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y119_SLICE_X27Y119_DO5),
.Q(\counter [17]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y119_SLICE_X27Y119_CARRY4 (
.CI(\$abc$3581$techmap2147$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[4].genblk1.carry4.genblk2.genblk1.cin_from_below ),
.CO({\$abc$3581$techmap2148$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[5].genblk1.carry4.genblk2.genblk1.cin_from_below , CLBLL_R_X17Y119_SLICE_X27Y119_C_CY, CLBLL_R_X17Y119_SLICE_X27Y119_B_CY, CLBLL_R_X17Y119_SLICE_X27Y119_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1415.Y [19], \$auto$alumacc.cc:485:replace_alu$1415.Y [18], \$auto$alumacc.cc:485:replace_alu$1415.Y [17], CLBLL_R_X17Y119_SLICE_X27Y119_A_XOR}),
.S({CLBLL_R_X17Y119_SLICE_X27Y119_DO6, CLBLL_R_X17Y119_SLICE_X27Y119_CO6, CLBLL_R_X17Y119_SLICE_X27Y119_BO6, CLBLL_R_X17Y119_SLICE_X27Y119_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLL_R_X17Y119_SLICE_X27Y119_DLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1415.Y [17]),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(\counter [19]),
.I5(1'b1),
.O5(CLBLL_R_X17Y119_SLICE_X27Y119_DO5),
.O6(CLBLL_R_X17Y119_SLICE_X27Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_R_X17Y119_SLICE_X27Y119_CLUT (
.I0(1'b1),
.I1(\$auto$alumacc.cc:485:replace_alu$1415.Y [19]),
.I2(\counter [18]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y119_SLICE_X27Y119_CO5),
.O6(CLBLL_R_X17Y119_SLICE_X27Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y119_SLICE_X27Y119_BLUT (
.I0(1'b1),
.I1(\counter [17]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1415.Y [18]),
.I5(1'b1),
.O5(CLBLL_R_X17Y119_SLICE_X27Y119_BO5),
.O6(CLBLL_R_X17Y119_SLICE_X27Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLL_R_X17Y119_SLICE_X27Y119_ALUT (
.I0(1'b1),
.I1(\counter [16]),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y119_SLICE_X27Y119_AO5),
.O6(CLBLL_R_X17Y119_SLICE_X27Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y120_SLICE_X26Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X26Y120_DO5),
.O6(CLBLL_R_X17Y120_SLICE_X26Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y120_SLICE_X26Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X26Y120_CO5),
.O6(CLBLL_R_X17Y120_SLICE_X26Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y120_SLICE_X26Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X26Y120_BO5),
.O6(CLBLL_R_X17Y120_SLICE_X26Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y120_SLICE_X26Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X26Y120_AO5),
.O6(CLBLL_R_X17Y120_SLICE_X26Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1523CLBLL_R_X17Y120_SLICE_X27Y120_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y120_SLICE_X27Y120_A_XOR),
.Q(\counter [20]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1525CLBLL_R_X17Y120_SLICE_X27Y120_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y120_SLICE_X27Y120_BO5),
.Q(\counter [22]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1526CLBLL_R_X17Y120_SLICE_X27Y120_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y120_SLICE_X27Y120_CO5),
.Q(\counter [23]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1524CLBLL_R_X17Y120_SLICE_X27Y120_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y120_SLICE_X27Y120_DO5),
.Q(\counter [21]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y120_SLICE_X27Y120_CARRY4 (
.CI(\$abc$3581$techmap2148$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[5].genblk1.carry4.genblk2.genblk1.cin_from_below ),
.CO({\$abc$3581$techmap2149$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[6].genblk1.carry4.genblk2.genblk1.cin_from_below , CLBLL_R_X17Y120_SLICE_X27Y120_C_CY, CLBLL_R_X17Y120_SLICE_X27Y120_B_CY, CLBLL_R_X17Y120_SLICE_X27Y120_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1415.Y [23], \$auto$alumacc.cc:485:replace_alu$1415.Y [22], \$auto$alumacc.cc:485:replace_alu$1415.Y [21], CLBLL_R_X17Y120_SLICE_X27Y120_A_XOR}),
.S({CLBLL_R_X17Y120_SLICE_X27Y120_DO6, CLBLL_R_X17Y120_SLICE_X27Y120_CO6, CLBLL_R_X17Y120_SLICE_X27Y120_BO6, CLBLL_R_X17Y120_SLICE_X27Y120_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_DLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1415.Y [21]),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(\counter [23]),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X27Y120_DO5),
.O6(CLBLL_R_X17Y120_SLICE_X27Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_CLUT (
.I0(1'b1),
.I1(\$auto$alumacc.cc:485:replace_alu$1415.Y [23]),
.I2(\counter [22]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X27Y120_CO5),
.O6(CLBLL_R_X17Y120_SLICE_X27Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_BLUT (
.I0(1'b1),
.I1(\counter [21]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1415.Y [22]),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X27Y120_BO5),
.O6(CLBLL_R_X17Y120_SLICE_X27Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLL_R_X17Y120_SLICE_X27Y120_ALUT (
.I0(1'b1),
.I1(\counter [20]),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y120_SLICE_X27Y120_AO5),
.O6(CLBLL_R_X17Y120_SLICE_X27Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y121_SLICE_X26Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y121_SLICE_X26Y121_DO5),
.O6(CLBLL_R_X17Y121_SLICE_X26Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y121_SLICE_X26Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y121_SLICE_X26Y121_CO5),
.O6(CLBLL_R_X17Y121_SLICE_X26Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y121_SLICE_X26Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y121_SLICE_X26Y121_BO5),
.O6(CLBLL_R_X17Y121_SLICE_X26Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y121_SLICE_X26Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y121_SLICE_X26Y121_AO5),
.O6(CLBLL_R_X17Y121_SLICE_X26Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1527CLBLL_R_X17Y121_SLICE_X27Y121_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y121_SLICE_X27Y121_A_XOR),
.Q(\counter [24]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1529CLBLL_R_X17Y121_SLICE_X27Y121_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y121_SLICE_X27Y121_BO5),
.Q(\counter [26]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1530CLBLL_R_X17Y121_SLICE_X27Y121_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y121_SLICE_X27Y121_CO5),
.Q(\counter [27]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:420:simplemap_dff$1528CLBLL_R_X17Y121_SLICE_X27Y121_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y121_SLICE_X27Y121_DO5),
.Q(\counter [25]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y121_SLICE_X27Y121_CARRY4 (
.CI(\$abc$3581$techmap2149$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[6].genblk1.carry4.genblk2.genblk1.cin_from_below ),
.CO({\$abc$3581$techmap2150$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[7].genblk1.carry4.genblk2.genblk1.cin_from_below , CLBLL_R_X17Y121_SLICE_X27Y121_C_CY, CLBLL_R_X17Y121_SLICE_X27Y121_B_CY, CLBLL_R_X17Y121_SLICE_X27Y121_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1415.Y [27], \$auto$alumacc.cc:485:replace_alu$1415.Y [26], \$auto$alumacc.cc:485:replace_alu$1415.Y [25], CLBLL_R_X17Y121_SLICE_X27Y121_A_XOR}),
.S({CLBLL_R_X17Y121_SLICE_X27Y121_DO6, CLBLL_R_X17Y121_SLICE_X27Y121_CO6, CLBLL_R_X17Y121_SLICE_X27Y121_BO6, CLBLL_R_X17Y121_SLICE_X27Y121_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLL_R_X17Y121_SLICE_X27Y121_DLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1415.Y [25]),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(\counter [27]),
.I5(1'b1),
.O5(CLBLL_R_X17Y121_SLICE_X27Y121_DO5),
.O6(CLBLL_R_X17Y121_SLICE_X27Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_R_X17Y121_SLICE_X27Y121_CLUT (
.I0(1'b1),
.I1(\$auto$alumacc.cc:485:replace_alu$1415.Y [27]),
.I2(\counter [26]),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y121_SLICE_X27Y121_CO5),
.O6(CLBLL_R_X17Y121_SLICE_X27Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_R_X17Y121_SLICE_X27Y121_BLUT (
.I0(1'b1),
.I1(\counter [25]),
.I2(1'b1),
.I3(1'b1),
.I4(\$auto$alumacc.cc:485:replace_alu$1415.Y [26]),
.I5(1'b1),
.O5(CLBLL_R_X17Y121_SLICE_X27Y121_BO5),
.O6(CLBLL_R_X17Y121_SLICE_X27Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLL_R_X17Y121_SLICE_X27Y121_ALUT (
.I0(1'b1),
.I1(\counter [24]),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y121_SLICE_X27Y121_AO5),
.O6(CLBLL_R_X17Y121_SLICE_X27Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y122_SLICE_X26Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y122_SLICE_X26Y122_DO5),
.O6(CLBLL_R_X17Y122_SLICE_X26Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y122_SLICE_X26Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y122_SLICE_X26Y122_CO5),
.O6(CLBLL_R_X17Y122_SLICE_X26Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y122_SLICE_X26Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y122_SLICE_X26Y122_BO5),
.O6(CLBLL_R_X17Y122_SLICE_X26Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y122_SLICE_X26Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y122_SLICE_X26Y122_AO5),
.O6(CLBLL_R_X17Y122_SLICE_X26Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y122_SLICE_X27Y122_A_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y122_SLICE_X27Y122_A_XOR),
.Q(CLBLL_R_X17Y122_SLICE_X27Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y122_SLICE_X27Y122_B_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y122_SLICE_X27Y122_BO5),
.Q(CLBLL_R_X17Y122_SLICE_X27Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y122_SLICE_X27Y122_C_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y122_SLICE_X27Y122_CO5),
.Q(CLBLL_R_X17Y122_SLICE_X27Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y122_SLICE_X27Y122_D_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y122_SLICE_X27Y122_DO5),
.Q(CLBLL_R_X17Y122_SLICE_X27Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y122_SLICE_X27Y122_CARRY4 (
.CI(\$abc$3581$techmap2150$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[7].genblk1.carry4.genblk2.genblk1.cin_from_below ),
.CO({\$abc$3581$techmap2151$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[8].genblk1.carry4.genblk2.genblk1.cin_from_below , CLBLL_R_X17Y122_SLICE_X27Y122_C_CY, CLBLL_R_X17Y122_SLICE_X27Y122_B_CY, CLBLL_R_X17Y122_SLICE_X27Y122_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1415.Y [31], \$auto$alumacc.cc:485:replace_alu$1415.Y [30], \$auto$alumacc.cc:485:replace_alu$1415.Y [29], CLBLL_R_X17Y122_SLICE_X27Y122_A_XOR}),
.S({CLBLL_R_X17Y122_SLICE_X27Y122_DO6, CLBLL_R_X17Y122_SLICE_X27Y122_CO6, CLBLL_R_X17Y122_SLICE_X27Y122_BO6, CLBLL_R_X17Y122_SLICE_X27Y122_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ff00)
  ) CLBLL_R_X17Y122_SLICE_X27Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_R_X17Y122_SLICE_X27Y122_CQ),
.I3(\$auto$alumacc.cc:485:replace_alu$1415.Y [29]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y122_SLICE_X27Y122_DO5),
.O6(CLBLL_R_X17Y122_SLICE_X27Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLL_R_X17Y122_SLICE_X27Y122_CLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1415.Y [31]),
.I1(CLBLL_R_X17Y122_SLICE_X27Y122_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y122_SLICE_X27Y122_CO5),
.O6(CLBLL_R_X17Y122_SLICE_X27Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLL_R_X17Y122_SLICE_X27Y122_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X17Y122_SLICE_X27Y122_DQ),
.I2(1'b1),
.I3(\$auto$alumacc.cc:485:replace_alu$1415.Y [30]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y122_SLICE_X27Y122_BO5),
.O6(CLBLL_R_X17Y122_SLICE_X27Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLL_R_X17Y122_SLICE_X27Y122_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X17Y122_SLICE_X27Y122_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y122_SLICE_X27Y122_AO5),
.O6(CLBLL_R_X17Y122_SLICE_X27Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y123_SLICE_X26Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y123_SLICE_X26Y123_DO5),
.O6(CLBLL_R_X17Y123_SLICE_X26Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y123_SLICE_X26Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y123_SLICE_X26Y123_CO5),
.O6(CLBLL_R_X17Y123_SLICE_X26Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y123_SLICE_X26Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y123_SLICE_X26Y123_BO5),
.O6(CLBLL_R_X17Y123_SLICE_X26Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X17Y123_SLICE_X26Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y123_SLICE_X26Y123_AO5),
.O6(CLBLL_R_X17Y123_SLICE_X26Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y123_SLICE_X27Y123_A_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y123_SLICE_X27Y123_A_XOR),
.Q(CLBLL_R_X17Y123_SLICE_X27Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y123_SLICE_X27Y123_B_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y123_SLICE_X27Y123_BO5),
.Q(CLBLL_R_X17Y123_SLICE_X27Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y123_SLICE_X27Y123_C_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y123_SLICE_X27Y123_CO5),
.Q(CLBLL_R_X17Y123_SLICE_X27Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X17Y123_SLICE_X27Y123_D_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLL_R_X17Y123_SLICE_X27Y123_DO5),
.Q(CLBLL_R_X17Y123_SLICE_X27Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_R_X17Y123_SLICE_X27Y123_CARRY4 (
.CI(\$abc$3581$techmap2151$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[8].genblk1.carry4.genblk2.genblk1.cin_from_below ),
.CO({CLBLL_R_X17Y123_SLICE_X27Y123_D_CY, CLBLL_R_X17Y123_SLICE_X27Y123_C_CY, CLBLL_R_X17Y123_SLICE_X27Y123_B_CY, CLBLL_R_X17Y123_SLICE_X27Y123_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({\$auto$alumacc.cc:485:replace_alu$1415.Y [35], \$auto$alumacc.cc:485:replace_alu$1415.Y [34], \$auto$alumacc.cc:485:replace_alu$1415.Y [33], CLBLL_R_X17Y123_SLICE_X27Y123_A_XOR}),
.S({CLBLL_R_X17Y123_SLICE_X27Y123_DO6, CLBLL_R_X17Y123_SLICE_X27Y123_CO6, CLBLL_R_X17Y123_SLICE_X27Y123_BO6, CLBLL_R_X17Y123_SLICE_X27Y123_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ff00)
  ) CLBLL_R_X17Y123_SLICE_X27Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_R_X17Y123_SLICE_X27Y123_CQ),
.I3(\$auto$alumacc.cc:485:replace_alu$1415.Y [33]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y123_SLICE_X27Y123_DO5),
.O6(CLBLL_R_X17Y123_SLICE_X27Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLL_R_X17Y123_SLICE_X27Y123_CLUT (
.I0(\$auto$alumacc.cc:485:replace_alu$1415.Y [35]),
.I1(CLBLL_R_X17Y123_SLICE_X27Y123_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y123_SLICE_X27Y123_CO5),
.O6(CLBLL_R_X17Y123_SLICE_X27Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLL_R_X17Y123_SLICE_X27Y123_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X17Y123_SLICE_X27Y123_DQ),
.I2(1'b1),
.I3(\$auto$alumacc.cc:485:replace_alu$1415.Y [34]),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y123_SLICE_X27Y123_BO5),
.O6(CLBLL_R_X17Y123_SLICE_X27Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLL_R_X17Y123_SLICE_X27Y123_ALUT (
.I0(1'b1),
.I1(CLBLL_R_X17Y123_SLICE_X27Y123_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X17Y123_SLICE_X27Y123_AO5),
.O6(CLBLL_R_X17Y123_SLICE_X27Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X43Y75_IOB_X1Y76_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O),
.O(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y1_OBUF (
.I(CLBLL_R_X17Y123_SLICE_X27Y123_CQ),
.O(led[7])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y2_OBUF (
.I(CLBLL_R_X17Y123_SLICE_X27Y123_BQ),
.O(led[6])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y121_IOB_X0Y122_IBUF (
.I(sw[3]),
.O(LIOB33_X0Y121_IOB_X0Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y123_IOB_X0Y123_IBUF (
.I(sw[2]),
.O(LIOB33_X0Y123_IOB_X0Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y123_IOB_X0Y124_IBUF (
.I(sw[1]),
.O(LIOB33_X0Y123_IOB_X0Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y125_IOB_X0Y125_IBUF (
.I(sw[0]),
.O(LIOB33_X0Y125_IOB_X0Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y125_IOB_X0Y126_IBUF (
.I(sw[7]),
.O(LIOB33_X0Y125_IOB_X0Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y127_IOB_X0Y127_IBUF (
.I(sw[6]),
.O(LIOB33_X0Y127_IOB_X0Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(sw[5]),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y137_IOB_X0Y137_IBUF (
.I(sw[4]),
.O(LIOB33_X0Y137_IOB_X0Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y51_IOB_X1Y51_OBUF (
.I(CLBLL_R_X17Y123_SLICE_X27Y123_AQ),
.O(led[4])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y51_IOB_X1Y52_OBUF (
.I(CLBLL_R_X17Y122_SLICE_X27Y122_CQ),
.O(led[3])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y55_IOB_X1Y55_OBUF (
.I(CLBLL_R_X17Y122_SLICE_X27Y122_BQ),
.O(led[2])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y57_IOB_X1Y58_OBUF (
.I(CLBLL_R_X17Y122_SLICE_X27Y122_DQ),
.O(led[1])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y61_IOB_X1Y61_OBUF (
.I(CLBLL_R_X17Y122_SLICE_X27Y122_AQ),
.O(led[0])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y75_IOB_X1Y76_IBUF (
.I(clk),
.O(RIOB33_X43Y75_IOB_X1Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_SING_X43Y50_IOB_X1Y50_OBUF (
.I(CLBLL_R_X17Y123_SLICE_X27Y123_DQ),
.O(led[5])
  );
  assign CLBLL_R_X17Y115_SLICE_X27Y115_COUT = \$abc$3581$techmap2144$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[1].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_AQ = \counter [0];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_BQ = \counter [2];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_CQ = \counter [3];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_DQ = \counter [1];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_BMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [1];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_CMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [2];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_DMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [3];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_COUT = \$abc$3581$techmap2145$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[2].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_AQ = \counter [6];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_BQ = \counter [7];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_CQ = \counter [4];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_DQ = \counter [5];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_AMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [4];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_BMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [5];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_CMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [6];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_DMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [7];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_COUT = \$abc$3581$techmap2146$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[3].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_AQ = \counter [10];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_BQ = \counter [11];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_CQ = \counter [8];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_DQ = \counter [9];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_AMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [8];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_BMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [9];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_CMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [10];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_DMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [11];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_COUT = \$abc$3581$techmap2147$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[4].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_AQ = \counter [14];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_BQ = \counter [15];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_CQ = \counter [12];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_DQ = \counter [13];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_AMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [12];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_BMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [13];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_CMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [14];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_DMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [15];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_COUT = \$abc$3581$techmap2148$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[5].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_AQ = \counter [16];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_BQ = \counter [18];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_CQ = \counter [19];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_DQ = \counter [17];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_BMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [17];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_CMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [18];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_DMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [19];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_COUT = \$abc$3581$techmap2149$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[6].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_AQ = \counter [20];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_BQ = \counter [22];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_CQ = \counter [23];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_DQ = \counter [21];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_BMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [21];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_CMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [22];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_DMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [23];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_COUT = \$abc$3581$techmap2150$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[7].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_AQ = \counter [24];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_BQ = \counter [26];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_CQ = \counter [27];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_DQ = \counter [25];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_BMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [25];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_CMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [26];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_DMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [27];
  assign CLBLL_R_X17Y122_SLICE_X27Y122_COUT = \$abc$3581$techmap2151$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[8].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_BMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [29];
  assign CLBLL_R_X17Y122_SLICE_X27Y122_CMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [30];
  assign CLBLL_R_X17Y122_SLICE_X27Y122_DMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [31];
  assign CLBLL_R_X17Y123_SLICE_X27Y123_BMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [33];
  assign CLBLL_R_X17Y123_SLICE_X27Y123_CMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [34];
  assign CLBLL_R_X17Y123_SLICE_X27Y123_DMUX = \$auto$alumacc.cc:485:replace_alu$1415.Y [35];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_B_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [1];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_C_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [2];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_D_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [3];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_D_CY = \$abc$3581$techmap2144$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[1].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_A_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [4];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_B_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [5];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_C_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [6];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_D_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [7];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_D_CY = \$abc$3581$techmap2145$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[2].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_A_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [8];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_B_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [9];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_C_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [10];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_D_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [11];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_D_CY = \$abc$3581$techmap2146$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[3].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_A_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [12];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_B_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [13];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_C_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [14];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [15];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D_CY = \$abc$3581$techmap2147$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[4].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_B_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [17];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_C_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [18];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [19];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D_CY = \$abc$3581$techmap2148$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[5].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [21];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [22];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [23];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D_CY = \$abc$3581$techmap2149$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[6].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_B_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [25];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_C_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [26];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [27];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D_CY = \$abc$3581$techmap2150$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[7].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_B_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [29];
  assign CLBLL_R_X17Y122_SLICE_X27Y122_C_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [30];
  assign CLBLL_R_X17Y122_SLICE_X27Y122_D_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [31];
  assign CLBLL_R_X17Y122_SLICE_X27Y122_D_CY = \$abc$3581$techmap2151$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[8].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_B_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [33];
  assign CLBLL_R_X17Y123_SLICE_X27Y123_C_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [34];
  assign CLBLL_R_X17Y123_SLICE_X27Y123_D_XOR = \$auto$alumacc.cc:485:replace_alu$1415.Y [35];
  assign CLBLL_R_X17Y115_SLICE_X26Y115_A = CLBLL_R_X17Y115_SLICE_X26Y115_AO6;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_B = CLBLL_R_X17Y115_SLICE_X26Y115_BO6;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_C = CLBLL_R_X17Y115_SLICE_X26Y115_CO6;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_D = CLBLL_R_X17Y115_SLICE_X26Y115_DO6;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_A = CLBLL_R_X17Y115_SLICE_X27Y115_AO6;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_B = CLBLL_R_X17Y115_SLICE_X27Y115_BO6;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_C = CLBLL_R_X17Y115_SLICE_X27Y115_CO6;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_D = CLBLL_R_X17Y115_SLICE_X27Y115_DO6;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_A = CLBLL_R_X17Y116_SLICE_X26Y116_AO6;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_B = CLBLL_R_X17Y116_SLICE_X26Y116_BO6;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_C = CLBLL_R_X17Y116_SLICE_X26Y116_CO6;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_D = CLBLL_R_X17Y116_SLICE_X26Y116_DO6;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_A = CLBLL_R_X17Y116_SLICE_X27Y116_AO6;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_B = CLBLL_R_X17Y116_SLICE_X27Y116_BO6;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_C = CLBLL_R_X17Y116_SLICE_X27Y116_CO6;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_D = CLBLL_R_X17Y116_SLICE_X27Y116_DO6;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_A = CLBLL_R_X17Y117_SLICE_X26Y117_AO6;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_B = CLBLL_R_X17Y117_SLICE_X26Y117_BO6;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_C = CLBLL_R_X17Y117_SLICE_X26Y117_CO6;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_D = CLBLL_R_X17Y117_SLICE_X26Y117_DO6;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_A = CLBLL_R_X17Y117_SLICE_X27Y117_AO6;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_B = CLBLL_R_X17Y117_SLICE_X27Y117_BO6;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_C = CLBLL_R_X17Y117_SLICE_X27Y117_CO6;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_D = CLBLL_R_X17Y117_SLICE_X27Y117_DO6;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_A = CLBLL_R_X17Y118_SLICE_X26Y118_AO6;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_B = CLBLL_R_X17Y118_SLICE_X26Y118_BO6;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_C = CLBLL_R_X17Y118_SLICE_X26Y118_CO6;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_D = CLBLL_R_X17Y118_SLICE_X26Y118_DO6;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_A = CLBLL_R_X17Y118_SLICE_X27Y118_AO6;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_B = CLBLL_R_X17Y118_SLICE_X27Y118_BO6;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_C = CLBLL_R_X17Y118_SLICE_X27Y118_CO6;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D = CLBLL_R_X17Y118_SLICE_X27Y118_DO6;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_A = CLBLL_R_X17Y119_SLICE_X26Y119_AO6;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_B = CLBLL_R_X17Y119_SLICE_X26Y119_BO6;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_C = CLBLL_R_X17Y119_SLICE_X26Y119_CO6;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_D = CLBLL_R_X17Y119_SLICE_X26Y119_DO6;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_A = CLBLL_R_X17Y119_SLICE_X27Y119_AO6;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_B = CLBLL_R_X17Y119_SLICE_X27Y119_BO6;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_C = CLBLL_R_X17Y119_SLICE_X27Y119_CO6;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D = CLBLL_R_X17Y119_SLICE_X27Y119_DO6;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A = CLBLL_R_X17Y120_SLICE_X26Y120_AO6;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B = CLBLL_R_X17Y120_SLICE_X26Y120_BO6;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C = CLBLL_R_X17Y120_SLICE_X26Y120_CO6;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D = CLBLL_R_X17Y120_SLICE_X26Y120_DO6;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A = CLBLL_R_X17Y120_SLICE_X27Y120_AO6;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B = CLBLL_R_X17Y120_SLICE_X27Y120_BO6;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C = CLBLL_R_X17Y120_SLICE_X27Y120_CO6;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D = CLBLL_R_X17Y120_SLICE_X27Y120_DO6;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_A = CLBLL_R_X17Y121_SLICE_X26Y121_AO6;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_B = CLBLL_R_X17Y121_SLICE_X26Y121_BO6;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_C = CLBLL_R_X17Y121_SLICE_X26Y121_CO6;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_D = CLBLL_R_X17Y121_SLICE_X26Y121_DO6;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_A = CLBLL_R_X17Y121_SLICE_X27Y121_AO6;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_B = CLBLL_R_X17Y121_SLICE_X27Y121_BO6;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_C = CLBLL_R_X17Y121_SLICE_X27Y121_CO6;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D = CLBLL_R_X17Y121_SLICE_X27Y121_DO6;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_A = CLBLL_R_X17Y122_SLICE_X26Y122_AO6;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_B = CLBLL_R_X17Y122_SLICE_X26Y122_BO6;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_C = CLBLL_R_X17Y122_SLICE_X26Y122_CO6;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_D = CLBLL_R_X17Y122_SLICE_X26Y122_DO6;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_A = CLBLL_R_X17Y122_SLICE_X27Y122_AO6;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_B = CLBLL_R_X17Y122_SLICE_X27Y122_BO6;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_C = CLBLL_R_X17Y122_SLICE_X27Y122_CO6;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_D = CLBLL_R_X17Y122_SLICE_X27Y122_DO6;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_A = CLBLL_R_X17Y123_SLICE_X26Y123_AO6;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_B = CLBLL_R_X17Y123_SLICE_X26Y123_BO6;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_C = CLBLL_R_X17Y123_SLICE_X26Y123_CO6;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_D = CLBLL_R_X17Y123_SLICE_X26Y123_DO6;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_A = CLBLL_R_X17Y123_SLICE_X27Y123_AO6;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_B = CLBLL_R_X17Y123_SLICE_X27Y123_BO6;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_C = CLBLL_R_X17Y123_SLICE_X27Y123_CO6;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_D = CLBLL_R_X17Y123_SLICE_X27Y123_DO6;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_OQ = CLBLL_R_X17Y123_SLICE_X27Y123_BQ;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_TQ = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_OQ = CLBLL_R_X17Y123_SLICE_X27Y123_CQ;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_TQ = 1'b1;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_O = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_O = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_O = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_O = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_OQ = CLBLL_R_X17Y122_SLICE_X27Y122_CQ;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_TQ = 1'b1;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_OQ = CLBLL_R_X17Y123_SLICE_X27Y123_AQ;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_TQ = 1'b1;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_OQ = CLBLL_R_X17Y122_SLICE_X27Y122_BQ;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_TQ = 1'b1;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_OQ = CLBLL_R_X17Y122_SLICE_X27Y122_AQ;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_TQ = 1'b1;
  assign RIOI3_X43Y75_ILOGIC_X1Y76_O = RIOB33_X43Y75_IOB_X1Y76_I;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_OQ = CLBLL_R_X17Y123_SLICE_X27Y123_DQ;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_OQ = CLBLL_R_X17Y122_SLICE_X27Y122_DQ;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_TQ = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_D1 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_D2 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_D3 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_D4 = \$auto$alumacc.cc:485:replace_alu$1415.Y [1];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_D5 = \counter [3];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_D6 = 1'b1;
  assign CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_CE = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_DX = 1'b0;
  assign LIOB33_X0Y1_IOB_X0Y2_O = CLBLL_R_X17Y123_SLICE_X27Y123_BQ;
  assign LIOB33_X0Y1_IOB_X0Y1_O = CLBLL_R_X17Y123_SLICE_X27Y123_CQ;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_D = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_A1 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_A2 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_A3 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_A4 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_A5 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_A6 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_B1 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_B2 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_B3 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_B4 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_B5 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_B6 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_C1 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_C2 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_C3 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_C4 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_C5 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_C6 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_D1 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_D2 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_D3 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_D4 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_D5 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X26Y122_D6 = 1'b1;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_D = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_A1 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_A2 = CLBLL_R_X17Y122_SLICE_X27Y122_AQ;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_A3 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_A4 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_A5 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_A6 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_AX = 1'b0;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_B1 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_B2 = CLBLL_R_X17Y122_SLICE_X27Y122_DQ;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_B3 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_B4 = \$auto$alumacc.cc:485:replace_alu$1415.Y [30];
  assign CLBLL_R_X17Y122_SLICE_X27Y122_B5 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_B6 = 1'b1;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_D1 = CLBLL_R_X17Y122_SLICE_X27Y122_BQ;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_BX = 1'b0;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_C1 = \$auto$alumacc.cc:485:replace_alu$1415.Y [31];
  assign CLBLL_R_X17Y122_SLICE_X27Y122_C2 = CLBLL_R_X17Y122_SLICE_X27Y122_BQ;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_C3 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_C4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_A1 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_A2 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_A3 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_A4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_A5 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_A6 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_C5 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_C6 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_CIN = \$abc$3581$techmap2150$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[7].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_B1 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_B2 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_B3 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_B4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_B5 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_B6 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_CX = 1'b0;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_D1 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_DX = 1'b0;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_C1 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_C2 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_C3 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_C4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_C5 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_C6 = 1'b1;
  assign RIOB33_X43Y57_IOB_X1Y58_O = CLBLL_R_X17Y122_SLICE_X27Y122_DQ;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_D1 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_D2 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_D3 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_D4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_D5 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X26Y119_D6 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_A1 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_A2 = \counter [16];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_A3 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_A4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_A5 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_A6 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_CX = 1'b0;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_AX = 1'b0;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_B1 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_B2 = \counter [17];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_B3 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_B4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_B5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [18];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_B6 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D1 = \$auto$alumacc.cc:485:replace_alu$1415.Y [17];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D2 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_BX = 1'b0;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_C1 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_C2 = \$auto$alumacc.cc:485:replace_alu$1415.Y [19];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_C3 = \counter [18];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_C4 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_A1 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_A2 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_A3 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_A4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_A5 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_A6 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_C5 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_C6 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_CIN = \$abc$3581$techmap2147$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[4].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_B1 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_B2 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D3 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D4 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D5 = \counter [19];
  assign CLBLL_R_X17Y119_SLICE_X27Y119_D6 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_B3 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_B4 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_B5 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_B6 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_C1 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_C2 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_C3 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_C4 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_C5 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_C6 = 1'b1;
  assign CLBLL_R_X17Y119_SLICE_X27Y119_DX = 1'b0;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_D1 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_D2 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_D3 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_D4 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_D5 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X26Y116_D6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D3 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D4 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D5 = \counter [27];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D6 = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_D = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_A1 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_A2 = \counter [4];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_A3 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_A4 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_A5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [6];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_A6 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_AX = 1'b0;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_B1 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_B2 = \counter [5];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_B3 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_B4 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_B5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [7];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_B6 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_BX = 1'b0;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_C1 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_C2 = \$auto$alumacc.cc:485:replace_alu$1415.Y [4];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_C3 = \counter [6];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_C4 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_C5 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_C6 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_D3 = CLBLL_R_X17Y123_SLICE_X27Y123_CQ;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_CIN = \$abc$3581$techmap2144$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[1].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_D4 = \$auto$alumacc.cc:485:replace_alu$1415.Y [33];
  assign CLBLL_R_X17Y123_SLICE_X27Y123_D5 = 1'b1;
  assign RIOB33_X43Y51_IOB_X1Y51_O = CLBLL_R_X17Y123_SLICE_X27Y123_AQ;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_CX = 1'b0;
  assign RIOB33_X43Y51_IOB_X1Y52_O = CLBLL_R_X17Y122_SLICE_X27Y122_CQ;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_D1 = \$auto$alumacc.cc:485:replace_alu$1415.Y [5];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_D2 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_D3 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_D4 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_D5 = \counter [7];
  assign CLBLL_R_X17Y116_SLICE_X27Y116_D6 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_D6 = 1'b1;
  assign CLBLL_R_X17Y116_SLICE_X27Y116_DX = 1'b0;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_A1 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_A2 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_A3 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_A4 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_A5 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_A6 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_B1 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_B2 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_B3 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_B4 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_B5 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_B6 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_C1 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_C2 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_C3 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_C4 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_C5 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_C6 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE0 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_CE1 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE0 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_IGNORE1 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S0 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_D1 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_D2 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_D3 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_D4 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_D5 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X26Y123_D6 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_S1 = 1'b1;
  assign RIOB33_SING_X43Y50_IOB_X1Y50_O = CLBLL_R_X17Y123_SLICE_X27Y123_DQ;
  assign RIOI3_X43Y75_ILOGIC_X1Y76_D = RIOB33_X43Y75_IOB_X1Y76_I;
  assign CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_I = CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_O;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_A1 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_A2 = CLBLL_R_X17Y123_SLICE_X27Y123_AQ;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_A3 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_A4 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_A5 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_A6 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_AX = 1'b0;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_B1 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_B2 = CLBLL_R_X17Y123_SLICE_X27Y123_DQ;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_B3 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_B4 = \$auto$alumacc.cc:485:replace_alu$1415.Y [34];
  assign CLBLL_R_X17Y123_SLICE_X27Y123_B5 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_B6 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_BX = 1'b0;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_C1 = \$auto$alumacc.cc:485:replace_alu$1415.Y [35];
  assign CLBLL_R_X17Y123_SLICE_X27Y123_C2 = CLBLL_R_X17Y123_SLICE_X27Y123_BQ;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_C3 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_C4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A2 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_A6 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_C5 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_C6 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_CIN = \$abc$3581$techmap2151$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[8].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B2 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_B6 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_CX = 1'b0;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_D1 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_D2 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C2 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_C6 = 1'b1;
  assign CLBLL_R_X17Y123_SLICE_X27Y123_DX = 1'b0;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D2 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X26Y120_D6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A2 = \counter [20];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_A6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_AX = 1'b0;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B2 = \counter [21];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B3 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B4 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [22];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_B6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_BX = 1'b0;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C2 = \$auto$alumacc.cc:485:replace_alu$1415.Y [23];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C3 = \counter [22];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C4 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_A1 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_A2 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_A3 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_A4 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_A5 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_A6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_C6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_CIN = \$abc$3581$techmap2148$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[5].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_B1 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_B2 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_B3 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_B4 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_B5 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_B6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_CX = 1'b0;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D1 = \$auto$alumacc.cc:485:replace_alu$1415.Y [21];
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D2 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_C1 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_C2 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_C3 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_C4 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_C5 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_C6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_DX = 1'b0;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_D = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_D1 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_D2 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_D3 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_D4 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_D5 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X26Y117_D6 = 1'b1;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_D = LIOB33_X0Y125_IOB_X0Y125_I;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_D1 = CLBLL_R_X17Y122_SLICE_X27Y122_AQ;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_T1 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_A1 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_A2 = \counter [8];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_A3 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_A4 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_A5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [10];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_A6 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_AX = 1'b0;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_B1 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_B2 = \counter [9];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_B3 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_B4 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_B5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [11];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_B6 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_BX = 1'b0;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_C1 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_C2 = \$auto$alumacc.cc:485:replace_alu$1415.Y [8];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_C3 = \counter [10];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_C4 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_C5 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_C6 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_CIN = \$abc$3581$techmap2145$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[2].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_CX = 1'b0;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_D1 = \$auto$alumacc.cc:485:replace_alu$1415.Y [9];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_D2 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_D3 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_D4 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_D5 = \counter [11];
  assign CLBLL_R_X17Y117_SLICE_X27Y117_D6 = 1'b1;
  assign CLBLL_R_X17Y117_SLICE_X27Y117_DX = 1'b0;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_D1 = CLBLL_R_X17Y122_SLICE_X27Y122_CQ;
  assign RIOI3_X43Y51_OLOGIC_X1Y52_T1 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_D1 = CLBLL_R_X17Y123_SLICE_X27Y123_BQ;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_D1 = CLBLL_R_X17Y123_SLICE_X27Y123_AQ;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_T1 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_CX = 1'b0;
  assign RIOI3_X43Y51_OLOGIC_X1Y51_T1 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_D1 = CLBLL_R_X17Y123_SLICE_X27Y123_CQ;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D1 = \$auto$alumacc.cc:485:replace_alu$1415.Y [13];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D2 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_T1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign RIOB33_X43Y61_IOB_X1Y61_O = CLBLL_R_X17Y122_SLICE_X27Y122_AQ;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_A1 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_A2 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_A3 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_A4 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_A5 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_A6 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D3 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_B1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D4 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_B2 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_B3 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_B4 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_B5 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D5 = \counter [23];
  assign CLBLL_R_X17Y121_SLICE_X26Y121_B6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_C1 = 1'b1;
  assign CLBLL_R_X17Y120_SLICE_X27Y120_D6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_C2 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_C3 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_C4 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_C5 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_D1 = CLBLL_R_X17Y122_SLICE_X27Y122_DQ;
  assign RIOI3_TBYTESRC_X43Y57_OLOGIC_X1Y58_T1 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_D1 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_D2 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_D3 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_D4 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_D5 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X26Y121_D6 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_D2 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_D3 = CLBLL_R_X17Y122_SLICE_X27Y122_CQ;
  assign RIOI3_X43Y55_OLOGIC_X1Y55_T1 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_D4 = \$auto$alumacc.cc:485:replace_alu$1415.Y [29];
  assign CLBLL_R_X17Y122_SLICE_X27Y122_D5 = 1'b1;
  assign CLBLL_R_X17Y122_SLICE_X27Y122_D6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_A1 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_A2 = \counter [24];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_A3 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_A4 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_A5 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_A6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_AX = 1'b0;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_B1 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_B2 = \counter [25];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_B3 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_B4 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_B5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [26];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_B6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_BX = 1'b0;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_C1 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_C2 = \$auto$alumacc.cc:485:replace_alu$1415.Y [27];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_C3 = \counter [26];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_C4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_A1 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_A2 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_A3 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_A4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_A5 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_A6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_C5 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_C6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_CIN = \$abc$3581$techmap2149$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[6].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_B1 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_B2 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_B3 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_B4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_B5 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_B6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_CX = 1'b0;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D1 = \$auto$alumacc.cc:485:replace_alu$1415.Y [25];
  assign CLBLL_R_X17Y121_SLICE_X27Y121_D2 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_C1 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_C2 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_C3 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_C4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_C5 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_C6 = 1'b1;
  assign CLBLL_R_X17Y121_SLICE_X27Y121_DX = 1'b0;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_D1 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_D2 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_D3 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_D4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_D5 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X26Y118_D6 = 1'b1;
  assign RIOB33_X43Y55_IOB_X1Y55_O = CLBLL_R_X17Y122_SLICE_X27Y122_BQ;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_D1 = CLBLL_R_X17Y123_SLICE_X27Y123_DQ;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_A1 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_A2 = \counter [12];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_A3 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_A4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_A5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [14];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_A6 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_AX = 1'b0;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_B1 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_B2 = \counter [13];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_B3 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_B4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_B5 = \$auto$alumacc.cc:485:replace_alu$1415.Y [15];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_B6 = 1'b1;
  assign RIOI3_SING_X43Y50_OLOGIC_X1Y50_T1 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_BX = 1'b0;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_C1 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_C2 = \$auto$alumacc.cc:485:replace_alu$1415.Y [12];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_C3 = \counter [14];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_C4 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_A1 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_A2 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_A3 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_A4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_A5 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_A6 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_C5 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_C6 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_CIN = \$abc$3581$techmap2146$auto$alumacc.cc:485:replace_alu$1415.genblk1.slice[3].genblk1.carry4.genblk2.genblk1.cin_from_below ;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_B1 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_B2 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D3 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D4 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D5 = \counter [15];
  assign CLBLL_R_X17Y118_SLICE_X27Y118_D6 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_B3 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_B4 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_B5 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_B6 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_C1 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_C2 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_C3 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_C4 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_C5 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_C6 = 1'b1;
  assign CLBLL_R_X17Y118_SLICE_X27Y118_DX = 1'b0;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_D1 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_D2 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_D3 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_D4 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_D5 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X26Y115_D6 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_A1 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_A2 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_A3 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_A4 = \counter [0];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_A5 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_A6 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_AX = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_B1 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_B2 = \counter [1];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_B3 = \$auto$alumacc.cc:485:replace_alu$1415.Y [2];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_B4 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_B5 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_B6 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_BX = 1'b0;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_C1 = \$auto$alumacc.cc:485:replace_alu$1415.Y [3];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_C2 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_C3 = \counter [2];
  assign CLBLL_R_X17Y115_SLICE_X27Y115_C4 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_C5 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_C6 = 1'b1;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I0 = RIOB33_X43Y75_IOB_X1Y76_I;
  assign CLK_BUFG_TOP_R_X60Y53_BUFGCTRL_X0Y16_I1 = 1'b1;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_D = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_R_X17Y115_SLICE_X27Y115_CX = 1'b0;
endmodule
