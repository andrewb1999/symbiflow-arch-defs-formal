module top(
  input clk,
  input rx,
  input [15:0] sw,
  output [15:0] led,
  output tx
  );
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR0;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR1;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR10;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR11;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR12;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR13;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR2;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR3;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR4;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR5;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR6;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR7;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR8;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR9;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRATIEHIGH0;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRATIEHIGH1;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBTIEHIGH0;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBTIEHIGH1;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR0;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR1;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR10;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR11;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR12;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR13;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR2;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR3;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR4;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR5;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR6;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR7;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR8;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR9;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIADI0;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIADI1;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIADI10;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIADI11;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIADI12;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIADI13;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIADI14;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIADI15;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIADI2;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIADI3;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIADI4;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIADI5;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIADI6;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIADI7;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIADI8;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIADI9;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI0;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI1;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI10;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI11;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI12;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI13;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI14;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI15;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI2;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI3;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI4;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI5;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI6;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI7;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI8;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI9;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIPADIP0;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIPADIP1;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIPBDIP0;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DIPBDIP1;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO0;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO1;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO10;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO11;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO12;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO13;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO14;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO15;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO16;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO17;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO18;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO19;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO2;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO20;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO21;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO22;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO23;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO24;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO25;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO26;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO27;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO28;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO29;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO3;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO30;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO31;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO4;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO5;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO6;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO7;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO8;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DO9;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DOP0;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DOP1;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DOP2;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_DOP3;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_RDCLK;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_RDEN;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_RDRCLK;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_REGCE;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_REGCEB;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_REGCLKB;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_RST;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_RSTRAMB;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_RSTREG;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_RSTREGB;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_WEA0;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_WEA1;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_WEA2;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_WEA3;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_WEBWE0;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_WEBWE1;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_WEBWE2;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_WEBWE3;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_WEBWE4;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_WEBWE5;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_WEBWE6;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_WEBWE7;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_WRCLK;
  wire [0:0] BRAM_L_X6Y120_RAMB18_X0Y48_WREN;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CLK;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D5Q;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CLK;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D5Q;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C5Q;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CLK;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D5Q;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C5Q;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CE;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CLK;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D5Q;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D5Q;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A5Q;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B5Q;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C5Q;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CE;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D5Q;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C5Q;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CLK;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D5Q;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C5Q;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CLK;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D5Q;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CLK;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C5Q;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CLK;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D5Q;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C5Q;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CE;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CLK;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D5Q;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B5Q;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C5Q;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CE;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CLK;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D5Q;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CE;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CLK;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_SR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_CE;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_I;
  wire [0:0] CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  wire [0:0] LIOB33_SING_X0Y0_IOB_X0Y0_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y11_I;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y12_I;
  wire [0:0] LIOB33_X0Y17_IOB_X0Y18_O;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y19_O;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y20_O;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_O;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y2_O;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y3_O;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y4_O;
  wire [0:0] LIOB33_X0Y43_IOB_X0Y43_O;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y5_I;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y6_I;
  wire [0:0] LIOB33_X0Y7_IOB_X0Y7_I;
  wire [0:0] LIOB33_X0Y7_IOB_X0Y8_I;
  wire [0:0] LIOB33_X0Y9_IOB_X0Y10_I;
  wire [0:0] LIOB33_X0Y9_IOB_X0Y9_I;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_D1;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_OQ;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_T1;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_O;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_O;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_D1;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_OQ;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_T1;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_TQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_TQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_TQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_D1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_OQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_T1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_TQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_D1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_OQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_T1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_TQ;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y5_D;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y5_O;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y6_D;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y6_O;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_D;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_O;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y9_D;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y9_O;
  wire [0:0] RIOB33_X43Y25_IOB_X1Y26_I;
  wire [0:0] RIOB33_X43Y31_IOB_X1Y32_O;
  wire [0:0] RIOB33_X43Y37_IOB_X1Y37_O;
  wire [0:0] RIOB33_X43Y37_IOB_X1Y38_O;
  wire [0:0] RIOB33_X43Y39_IOB_X1Y39_I;
  wire [0:0] RIOB33_X43Y39_IOB_X1Y40_I;
  wire [0:0] RIOB33_X43Y43_IOB_X1Y43_I;
  wire [0:0] RIOB33_X43Y43_IOB_X1Y44_I;
  wire [0:0] RIOB33_X43Y45_IOB_X1Y45_I;
  wire [0:0] RIOB33_X43Y45_IOB_X1Y46_I;
  wire [0:0] RIOB33_X43Y47_IOB_X1Y47_I;
  wire [0:0] RIOB33_X43Y47_IOB_X1Y48_I;
  wire [0:0] RIOB33_X43Y61_IOB_X1Y61_O;
  wire [0:0] RIOB33_X43Y75_IOB_X1Y75_O;
  wire [0:0] RIOB33_X43Y75_IOB_X1Y76_O;
  wire [0:0] RIOB33_X43Y87_IOB_X1Y87_O;
  wire [0:0] RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_D1;
  wire [0:0] RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_OQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_T1;
  wire [0:0] RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_TQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y43_D;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y43_O;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y44_D;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y44_O;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_D1;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_OQ;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_T1;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_TQ;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_D1;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_OQ;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_T1;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_TQ;
  wire [0:0] RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_D1;
  wire [0:0] RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_OQ;
  wire [0:0] RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_T1;
  wire [0:0] RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_TQ;
  wire [0:0] RIOI3_X43Y25_ILOGIC_X1Y26_D;
  wire [0:0] RIOI3_X43Y25_ILOGIC_X1Y26_O;
  wire [0:0] RIOI3_X43Y39_ILOGIC_X1Y39_D;
  wire [0:0] RIOI3_X43Y39_ILOGIC_X1Y39_O;
  wire [0:0] RIOI3_X43Y39_ILOGIC_X1Y40_D;
  wire [0:0] RIOI3_X43Y39_ILOGIC_X1Y40_O;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y45_D;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y45_O;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y46_D;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y46_O;
  wire [0:0] RIOI3_X43Y47_ILOGIC_X1Y47_D;
  wire [0:0] RIOI3_X43Y47_ILOGIC_X1Y47_O;
  wire [0:0] RIOI3_X43Y47_ILOGIC_X1Y48_D;
  wire [0:0] RIOI3_X43Y47_ILOGIC_X1Y48_O;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_D1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_OQ;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_T1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_TQ;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y75_D1;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y75_OQ;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y75_T1;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y75_TQ;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y76_D1;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y76_OQ;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y76_T1;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y76_TQ;
  wire [0:0] \$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1517 ;
  wire [0:0] \$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1522 ;
  wire [0:0] \$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1525 ;
  wire [0:0] \$abc$2590$auto$rtlil.cc:2282:AndGate$1870 ;
  wire [0:0] \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2657 ;
  wire [0:0] \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2659 ;
  wire [0:0] \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2661 ;
  wire [0:0] \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2663 ;
  wire [0:0] \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2665 ;
  wire [0:0] \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2667 ;
  wire [1:0] \$techmap2616$abc$2590$lut$auto$opt_dff.cc:242:make_patterns_logic$1522.A ;
  wire [15:0] \ram.di ;
  wire [15:0] \ram.do ;
  wire [9:0] \wraddr ;
  wire [0:0] \wren ;


  (* KEEP, DONT_TOUCH, BEL = "RAMB18E1" *)
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000004450),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000000040002193366CC070F78F07FFF2A5555AA0001),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .IS_CLKARDCLK_INVERTED(0),
    .IS_CLKBWRCLK_INVERTED(0),
    .IS_ENARDEN_INVERTED(0),
    .IS_ENBWREN_INVERTED(0),
    .IS_RSTRAMARSTRAM_INVERTED(1),
    .IS_RSTRAMB_INVERTED(1),
    .IS_RSTREGARSTREG_INVERTED(1),
    .IS_RSTREGB_INVERTED(1),
    .RAM_MODE("TDP"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("READ_FIRST"),
    .WRITE_MODE_B("READ_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(18)
  ) \ram.ram.0.0.0BRAM_L_X6Y120_RAMB18_X0Y48_RAMB18E1  (
.ADDRARDADDR({\wraddr [9], \wraddr [8], \wraddr [7], \wraddr [6], \wraddr [5], \wraddr [4], \wraddr [3], \wraddr [2], \wraddr [1], \wraddr [0], 1'b0, 1'b0, 1'b0, 1'b0}),
.ADDRBWRADDR({\wraddr [9], \wraddr [8], \wraddr [7], \wraddr [6], \wraddr [5], \wraddr [4], \wraddr [3], \wraddr [2], \wraddr [1], \wraddr [0], 1'b0, 1'b0, 1'b0, 1'b0}),
.CLKARDCLK(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CLKBWRCLK(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.DIADI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.DIBDI({1'b0, \ram.di [15], \ram.di [14], \ram.di [13], \ram.di [12], \ram.di [11], \ram.di [10], \ram.di [9], \ram.di [7], \ram.di [6], \ram.di [5], \ram.di [4], \ram.di [3], \ram.di [2], \ram.di [1], \ram.di [0]}),
.DIPADIP({1'b0, 1'b0}),
.DIPBDIP({1'b0, \ram.di [8]}),
.DOADO({BRAM_L_X6Y120_RAMB18_X0Y48_DO15, \ram.do [15], \ram.do [14], \ram.do [13], \ram.do [12], \ram.do [11], \ram.do [10], \ram.do [9], \ram.do [7], \ram.do [6], \ram.do [5], \ram.do [4], \ram.do [3], \ram.do [2], \ram.do [1], \ram.do [0]}),
.DOBDO({BRAM_L_X6Y120_RAMB18_X0Y48_DO31, BRAM_L_X6Y120_RAMB18_X0Y48_DO30, BRAM_L_X6Y120_RAMB18_X0Y48_DO29, BRAM_L_X6Y120_RAMB18_X0Y48_DO28, BRAM_L_X6Y120_RAMB18_X0Y48_DO27, BRAM_L_X6Y120_RAMB18_X0Y48_DO26, BRAM_L_X6Y120_RAMB18_X0Y48_DO25, BRAM_L_X6Y120_RAMB18_X0Y48_DO24, BRAM_L_X6Y120_RAMB18_X0Y48_DO23, BRAM_L_X6Y120_RAMB18_X0Y48_DO22, BRAM_L_X6Y120_RAMB18_X0Y48_DO21, BRAM_L_X6Y120_RAMB18_X0Y48_DO20, BRAM_L_X6Y120_RAMB18_X0Y48_DO19, BRAM_L_X6Y120_RAMB18_X0Y48_DO18, BRAM_L_X6Y120_RAMB18_X0Y48_DO17, BRAM_L_X6Y120_RAMB18_X0Y48_DO16}),
.DOPADOP({BRAM_L_X6Y120_RAMB18_X0Y48_DOP1, \ram.do [8]}),
.DOPBDOP({BRAM_L_X6Y120_RAMB18_X0Y48_DOP3, BRAM_L_X6Y120_RAMB18_X0Y48_DOP2}),
.ENARDEN(1'b1),
.ENBWREN(1'b1),
.REGCEAREGCE(1'b1),
.REGCEB(1'b0),
.RSTRAMARSTRAM(1'b1),
.RSTRAMB(1'b1),
.RSTREGARSTREG(1'b1),
.RSTREGB(1'b1),
.WEA({1'b0, 1'b0}),
.WEBWE({\wren , \wren })
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_C5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$abc$4086$auto$xilinx_dffopt.cc:347:execute$2663 ),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_D5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$abc$4086$auto$xilinx_dffopt.cc:347:execute$2661 ),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_DO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_CO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cf0ac00a)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_BLUT (
.I0(\ram.do [13]),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.I2(RIOB33_X43Y43_IOB_X1Y44_I),
.I3(RIOB33_X43Y47_IOB_X1Y48_I),
.I4(\ram.di [13]),
.I5(1'b1),
.O5(\$abc$4086$auto$xilinx_dffopt.cc:347:execute$2663 ),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cbc80b08)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_ALUT (
.I0(\ram.di [12]),
.I1(RIOB33_X43Y47_IOB_X1Y48_I),
.I2(RIOB33_X43Y43_IOB_X1Y44_I),
.I3(\ram.do [12]),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_D5Q),
.I5(1'b1),
.O5(\$abc$4086$auto$xilinx_dffopt.cc:347:execute$2661 ),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_C5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$abc$4086$auto$xilinx_dffopt.cc:347:execute$2667 ),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_D5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$abc$4086$auto$xilinx_dffopt.cc:347:execute$2657 ),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_DO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_CO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cf0ac00a)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_BLUT (
.I0(\ram.do [15]),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_C5Q),
.I2(RIOB33_X43Y43_IOB_X1Y44_I),
.I3(RIOB33_X43Y47_IOB_X1Y48_I),
.I4(\ram.di [15]),
.I5(1'b1),
.O5(\$abc$4086$auto$xilinx_dffopt.cc:347:execute$2667 ),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cbc80b08)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_ALUT (
.I0(\ram.di [10]),
.I1(RIOB33_X43Y47_IOB_X1Y48_I),
.I2(RIOB33_X43Y43_IOB_X1Y44_I),
.I3(\ram.do [10]),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_D5Q),
.I5(1'b1),
.O5(\$abc$4086$auto$xilinx_dffopt.cc:347:execute$2657 ),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_C5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_BO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_D5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_AO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfadd50ddfa885088)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_BLUT (
.I0(RIOB33_X43Y43_IOB_X1Y44_I),
.I1(\wraddr [7]),
.I2(\ram.di [7]),
.I3(RIOB33_X43Y47_IOB_X1Y48_I),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_C5Q),
.I5(\ram.do [7]),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefe32f23ece02c20)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_ALUT (
.I0(\ram.di [2]),
.I1(RIOB33_X43Y43_IOB_X1Y44_I),
.I2(RIOB33_X43Y47_IOB_X1Y48_I),
.I3(\wraddr [2]),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_D5Q),
.I5(\ram.do [2]),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1758CLBLM_R_X5Y119_SLICE_X7Y119_C5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1525 ),
.D(LIOB33_X0Y7_IOB_X0Y7_I),
.Q(\wraddr [4]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1755CLBLM_R_X5Y119_SLICE_X7Y119_D5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1525 ),
.D(LIOB33_X0Y11_IOB_X0Y12_I),
.Q(\wraddr [1]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1756CLBLM_R_X5Y119_SLICE_X7Y119_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1525 ),
.D(CLBLM_R_X5Y119_SLICE_X7Y119_CO5),
.Q(\wraddr [2]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1757CLBLM_R_X5Y119_SLICE_X7Y119_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1525 ),
.D(CLBLM_R_X5Y119_SLICE_X7Y119_DO5),
.Q(\wraddr [3]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y9_IOB_X0Y9_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff0000)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y9_IOB_X0Y10_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_C5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_BO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_D5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_AO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfadd50ddfa885088)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_BLUT (
.I0(RIOB33_X43Y43_IOB_X1Y44_I),
.I1(\wraddr [8]),
.I2(\ram.di [8]),
.I3(RIOB33_X43Y47_IOB_X1Y48_I),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_C5Q),
.I5(\ram.do [8]),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefe32f23ece02c20)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_ALUT (
.I0(\ram.di [1]),
.I1(RIOB33_X43Y43_IOB_X1Y44_I),
.I2(RIOB33_X43Y47_IOB_X1Y48_I),
.I3(\wraddr [1]),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_D5Q),
.I5(\ram.do [1]),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1767CLBLM_R_X5Y120_SLICE_X7Y120_A5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1522 ),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_AO5),
.Q(\ram.di [1]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1768CLBLM_R_X5Y120_SLICE_X7Y120_B5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1522 ),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_BO5),
.Q(\ram.di [2]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1773CLBLM_R_X5Y120_SLICE_X7Y120_C5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1522 ),
.D(LIOB33_X0Y5_IOB_X0Y6_I),
.Q(\ram.di [7]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1766CLBLM_R_X5Y120_SLICE_X7Y120_D5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1522 ),
.D(LIOB33_X0Y11_IOB_X0Y11_I),
.Q(\ram.di [0]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1769CLBLM_R_X5Y120_SLICE_X7Y120_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1522 ),
.D(LIOB33_X0Y9_IOB_X0Y9_I),
.Q(\ram.di [3]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1770CLBLM_R_X5Y120_SLICE_X7Y120_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1522 ),
.D(LIOB33_X0Y7_IOB_X0Y7_I),
.Q(\ram.di [4]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1771CLBLM_R_X5Y120_SLICE_X7Y120_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1522 ),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_CO5),
.Q(\ram.di [5]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1772CLBLM_R_X5Y120_SLICE_X7Y120_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1522 ),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_DO5),
.Q(\ram.di [6]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y5_IOB_X0Y5_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y7_IOB_X0Y8_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff0000)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y9_IOB_X0Y10_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y11_IOB_X0Y12_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_C5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_BO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_D5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_AO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_DO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_CO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfadd50ddfa885088)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_BLUT (
.I0(RIOB33_X43Y43_IOB_X1Y44_I),
.I1(\wraddr [6]),
.I2(\ram.di [6]),
.I3(RIOB33_X43Y47_IOB_X1Y48_I),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_C5Q),
.I5(\ram.do [6]),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_BO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbcb3b0bf8c83808)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_ALUT (
.I0(\wraddr [3]),
.I1(RIOB33_X43Y43_IOB_X1Y44_I),
.I2(RIOB33_X43Y47_IOB_X1Y48_I),
.I3(\ram.di [3]),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_D5Q),
.I5(\ram.do [3]),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_AO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_C5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X7Y121_BO6),
.Q(CLBLM_R_X5Y121_SLICE_X7Y121_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_D5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X7Y121_AO6),
.Q(CLBLM_R_X5Y121_SLICE_X7Y121_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_DO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_CO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfadd50ddfa885088)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_BLUT (
.I0(RIOB33_X43Y43_IOB_X1Y44_I),
.I1(\wraddr [5]),
.I2(\ram.di [5]),
.I3(RIOB33_X43Y47_IOB_X1Y48_I),
.I4(CLBLM_R_X5Y121_SLICE_X7Y121_C5Q),
.I5(\ram.do [5]),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_BO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefe32f23ece02c20)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_ALUT (
.I0(\ram.di [4]),
.I1(RIOB33_X43Y43_IOB_X1Y44_I),
.I2(RIOB33_X43Y47_IOB_X1Y48_I),
.I3(\wraddr [4]),
.I4(CLBLM_R_X5Y121_SLICE_X7Y121_D5Q),
.I5(\ram.do [4]),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_AO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_C5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_BO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_D5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_AO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heef544f5eea044a0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_BLUT (
.I0(RIOB33_X43Y43_IOB_X1Y44_I),
.I1(\ram.di [9]),
.I2(\wraddr [9]),
.I3(RIOB33_X43Y47_IOB_X1Y48_I),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_C5Q),
.I5(\ram.do [9]),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbcb3b0bf8c83808)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_ALUT (
.I0(\wraddr [0]),
.I1(RIOB33_X43Y43_IOB_X1Y44_I),
.I2(RIOB33_X43Y47_IOB_X1Y48_I),
.I3(\ram.di [0]),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_D5Q),
.I5(\ram.do [0]),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_C5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$abc$4086$auto$xilinx_dffopt.cc:347:execute$2665 ),
.Q(CLBLM_R_X7Y119_SLICE_X9Y119_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_D5_FDRE (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(1'b1),
.D(\$abc$4086$auto$xilinx_dffopt.cc:347:execute$2659 ),
.Q(CLBLM_R_X7Y119_SLICE_X9Y119_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cf0ac00a)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_BLUT (
.I0(\ram.do [14]),
.I1(CLBLM_R_X7Y119_SLICE_X9Y119_C5Q),
.I2(RIOB33_X43Y43_IOB_X1Y44_I),
.I3(RIOB33_X43Y47_IOB_X1Y48_I),
.I4(\ram.di [14]),
.I5(1'b1),
.O5(\$abc$4086$auto$xilinx_dffopt.cc:347:execute$2665 ),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cbc80b08)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_ALUT (
.I0(\ram.di [11]),
.I1(RIOB33_X43Y47_IOB_X1Y48_I),
.I2(RIOB33_X43Y43_IOB_X1Y44_I),
.I3(\ram.do [11]),
.I4(CLBLM_R_X7Y119_SLICE_X9Y119_D5Q),
.I5(1'b1),
.O5(\$abc$4086$auto$xilinx_dffopt.cc:347:execute$2659 ),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1763CLBLM_R_X7Y120_SLICE_X8Y120_C5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1525 ),
.D(RIOB33_X43Y45_IOB_X1Y45_I),
.Q(\wraddr [9]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1754CLBLM_R_X7Y120_SLICE_X8Y120_D5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1525 ),
.D(LIOB33_X0Y11_IOB_X0Y11_I),
.Q(\wraddr [0]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1759CLBLM_R_X7Y120_SLICE_X8Y120_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1525 ),
.D(LIOB33_X0Y7_IOB_X0Y8_I),
.Q(\wraddr [5]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1760CLBLM_R_X7Y120_SLICE_X8Y120_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1525 ),
.D(LIOB33_X0Y5_IOB_X0Y5_I),
.Q(\wraddr [6]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1761CLBLM_R_X7Y120_SLICE_X8Y120_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1525 ),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_CO5),
.Q(\wraddr [7]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1762CLBLM_R_X7Y120_SLICE_X8Y120_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1525 ),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_DO5),
.Q(\wraddr [8]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h20202020ffff0000)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_DLUT (
.I0(RIOB33_X43Y45_IOB_X1Y46_I),
.I1(RIOB33_X43Y39_IOB_X1Y39_I),
.I2(RIOB33_X43Y43_IOB_X1Y43_I),
.I3(1'b1),
.I4(RIOB33_X43Y39_IOB_X1Y40_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_DO5),
.O6(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1517 )
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y5_IOB_X0Y6_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2a2a2a2acccc0000)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_BLUT (
.I0(RIOB33_X43Y45_IOB_X1Y46_I),
.I1(RIOB33_X43Y39_IOB_X1Y39_I),
.I2(RIOB33_X43Y43_IOB_X1Y43_I),
.I3(1'b1),
.I4(\$techmap2616$abc$2590$lut$auto$opt_dff.cc:242:make_patterns_logic$1522.A [1]),
.I5(1'b1),
.O5(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1522 ),
.O6(\$abc$2590$auto$rtlil.cc:2282:AndGate$1870 )
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff0044444444)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_ALUT (
.I0(RIOB33_X43Y39_IOB_X1Y39_I),
.I1(\$techmap2616$abc$2590$lut$auto$opt_dff.cc:242:make_patterns_logic$1522.A [1]),
.I2(1'b1),
.I3(RIOB33_X43Y45_IOB_X1Y46_I),
.I4(RIOB33_X43Y43_IOB_X1Y43_I),
.I5(1'b1),
.O5(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1525 ),
.O6(\$techmap2616$abc$2590$lut$auto$opt_dff.cc:242:make_patterns_logic$1522.A [1])
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1677CLBLM_R_X7Y120_SLICE_X9Y120_A5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1517 ),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_AO5),
.Q(\ram.di [9]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1678CLBLM_R_X7Y120_SLICE_X9Y120_B5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1517 ),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_BO5),
.Q(\ram.di [10]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1683CLBLM_R_X7Y120_SLICE_X9Y120_C5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1517 ),
.D(LIOB33_X0Y5_IOB_X0Y6_I),
.Q(\ram.di [15]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1676CLBLM_R_X7Y120_SLICE_X9Y120_D5_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1517 ),
.D(LIOB33_X0Y11_IOB_X0Y11_I),
.Q(\ram.di [8]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1679CLBLM_R_X7Y120_SLICE_X9Y120_A_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1517 ),
.D(LIOB33_X0Y9_IOB_X0Y9_I),
.Q(\ram.di [11]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1680CLBLM_R_X7Y120_SLICE_X9Y120_B_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1517 ),
.D(LIOB33_X0Y7_IOB_X0Y7_I),
.Q(\ram.di [12]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1681CLBLM_R_X7Y120_SLICE_X9Y120_C_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1517 ),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_CO5),
.Q(\ram.di [13]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:442:simplemap_dffe$1682CLBLM_R_X7Y120_SLICE_X9Y120_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(\$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1517 ),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_DO5),
.Q(\ram.di [14]),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y5_IOB_X0Y5_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y7_IOB_X0Y8_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff0000)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y9_IOB_X0Y10_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y11_IOB_X0Y12_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) \$auto$simplemap.cc:559:simplemap_adffe_sdffe_sdffce$1726CLBLM_R_X7Y121_SLICE_X8Y121_D_FDRE  (
.C(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O),
.CE(RIOB33_X43Y45_IOB_X1Y46_I),
.D(1'b1),
.Q(\wren ),
.R(\$abc$2590$auto$rtlil.cc:2282:AndGate$1870 )
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X43Y25_IOB_X1Y26_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y1_OBUF (
.I(CLBLM_R_X5Y119_SLICE_X6Y119_C5Q),
.O(led[7])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y2_OBUF (
.I(CLBLM_R_X5Y120_SLICE_X6Y120_C5Q),
.O(led[8])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y3_IOB_X0Y3_OBUF (
.I(CLBLM_R_X7Y119_SLICE_X8Y119_D5Q),
.O(led[0])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y3_IOB_X0Y4_OBUF (
.I(CLBLM_R_X5Y121_SLICE_X7Y121_C5Q),
.O(led[5])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y5_IOB_X0Y5_IBUF (
.I(sw[6]),
.O(LIOB33_X0Y5_IOB_X0Y5_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y5_IOB_X0Y6_IBUF (
.I(sw[7]),
.O(LIOB33_X0Y5_IOB_X0Y6_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y7_IOB_X0Y7_IBUF (
.I(sw[4]),
.O(LIOB33_X0Y7_IOB_X0Y7_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y7_IOB_X0Y8_IBUF (
.I(sw[5]),
.O(LIOB33_X0Y7_IOB_X0Y8_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y9_IOB_X0Y9_IBUF (
.I(sw[3]),
.O(LIOB33_X0Y9_IOB_X0Y9_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y9_IOB_X0Y10_IBUF (
.I(sw[2]),
.O(LIOB33_X0Y9_IOB_X0Y10_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y11_IOB_X0Y11_IBUF (
.I(sw[0]),
.O(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y11_IOB_X0Y12_IBUF (
.I(sw[1]),
.O(LIOB33_X0Y11_IOB_X0Y12_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y17_IOB_X0Y18_OBUF (
.I(CLBLM_R_X5Y121_SLICE_X7Y121_D5Q),
.O(led[4])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y19_IOB_X0Y19_OBUF (
.I(CLBLM_R_X5Y121_SLICE_X6Y121_D5Q),
.O(led[3])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y19_IOB_X0Y20_OBUF (
.I(CLBLM_R_X5Y119_SLICE_X6Y119_D5Q),
.O(led[2])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y43_IOB_X0Y43_OBUF (
.I(CLBLM_R_X5Y120_SLICE_X6Y120_D5Q),
.O(led[1])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_I),
.O(tx)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(rx),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y0_IOB_X0Y0_OBUF (
.I(CLBLM_R_X5Y121_SLICE_X6Y121_C5Q),
.O(led[6])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y25_IOB_X1Y26_IBUF (
.I(clk),
.O(RIOB33_X43Y25_IOB_X1Y26_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y31_IOB_X1Y32_OBUF (
.I(CLBLM_R_X7Y119_SLICE_X9Y119_D5Q),
.O(led[11])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y37_IOB_X1Y37_OBUF (
.I(CLBLM_L_X8Y120_SLICE_X11Y120_D5Q),
.O(led[10])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y37_IOB_X1Y38_OBUF (
.I(CLBLM_R_X7Y119_SLICE_X8Y119_C5Q),
.O(led[9])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y39_IOB_X1Y39_IBUF (
.I(sw[12]),
.O(RIOB33_X43Y39_IOB_X1Y39_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y39_IOB_X1Y40_IBUF (
.I(sw[8]),
.O(RIOB33_X43Y39_IOB_X1Y40_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y43_IOB_X1Y43_IBUF (
.I(sw[13]),
.O(RIOB33_X43Y43_IOB_X1Y43_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y43_IOB_X1Y44_IBUF (
.I(sw[14]),
.O(RIOB33_X43Y43_IOB_X1Y44_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y45_IOB_X1Y45_IBUF (
.I(sw[9]),
.O(RIOB33_X43Y45_IOB_X1Y45_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y45_IOB_X1Y46_IBUF (
.I(sw[11]),
.O(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y47_IOB_X1Y47_IBUF (
.I(sw[10]),
.O(RIOB33_X43Y47_IOB_X1Y47_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y47_IOB_X1Y48_IBUF (
.I(sw[15]),
.O(RIOB33_X43Y47_IOB_X1Y48_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y61_IOB_X1Y61_OBUF (
.I(CLBLM_R_X7Y119_SLICE_X9Y119_C5Q),
.O(led[14])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y75_IOB_X1Y75_OBUF (
.I(CLBLM_L_X8Y120_SLICE_X10Y120_D5Q),
.O(led[12])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y75_IOB_X1Y76_OBUF (
.I(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.O(led[13])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y87_IOB_X1Y87_OBUF (
.I(CLBLM_L_X8Y120_SLICE_X11Y120_C5Q),
.O(led[15])
  );
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DO0 = \ram.do [0];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DO1 = \ram.do [1];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DO2 = \ram.do [2];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DO3 = \ram.do [3];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DO4 = \ram.do [4];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DO5 = \ram.do [5];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DO6 = \ram.do [6];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DO7 = \ram.do [7];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DO8 = \ram.do [9];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DO9 = \ram.do [10];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DO10 = \ram.do [11];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DO11 = \ram.do [12];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DO12 = \ram.do [13];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DO13 = \ram.do [14];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DO14 = \ram.do [15];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DOP0 = \ram.do [8];
  assign CLBLM_L_X8Y120_SLICE_X10Y120_AMUX = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2661 ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_BMUX = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2663 ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_AMUX = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2657 ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_BMUX = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2667 ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_CQ = \wraddr [2];
  assign CLBLM_R_X5Y119_SLICE_X7Y119_DQ = \wraddr [3];
  assign CLBLM_R_X5Y119_SLICE_X7Y119_CMUX = \wraddr [4];
  assign CLBLM_R_X5Y119_SLICE_X7Y119_DMUX = \wraddr [1];
  assign CLBLM_R_X5Y120_SLICE_X7Y120_AQ = \ram.di [3];
  assign CLBLM_R_X5Y120_SLICE_X7Y120_BQ = \ram.di [4];
  assign CLBLM_R_X5Y120_SLICE_X7Y120_CQ = \ram.di [5];
  assign CLBLM_R_X5Y120_SLICE_X7Y120_DQ = \ram.di [6];
  assign CLBLM_R_X5Y120_SLICE_X7Y120_AMUX = \ram.di [1];
  assign CLBLM_R_X5Y120_SLICE_X7Y120_BMUX = \ram.di [2];
  assign CLBLM_R_X5Y120_SLICE_X7Y120_CMUX = \ram.di [7];
  assign CLBLM_R_X5Y120_SLICE_X7Y120_DMUX = \ram.di [0];
  assign CLBLM_R_X7Y119_SLICE_X9Y119_AMUX = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2659 ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_BMUX = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2665 ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_AQ = \wraddr [5];
  assign CLBLM_R_X7Y120_SLICE_X8Y120_BQ = \wraddr [6];
  assign CLBLM_R_X7Y120_SLICE_X8Y120_CQ = \wraddr [7];
  assign CLBLM_R_X7Y120_SLICE_X8Y120_DQ = \wraddr [8];
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A = \$techmap2616$abc$2590$lut$auto$opt_dff.cc:242:make_patterns_logic$1522.A [1];
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B = \$abc$2590$auto$rtlil.cc:2282:AndGate$1870 ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D = \$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1517 ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_AMUX = \$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1525 ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_BMUX = \$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1522 ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_CMUX = \wraddr [9];
  assign CLBLM_R_X7Y120_SLICE_X8Y120_DMUX = \wraddr [0];
  assign CLBLM_R_X7Y120_SLICE_X9Y120_AQ = \ram.di [11];
  assign CLBLM_R_X7Y120_SLICE_X9Y120_BQ = \ram.di [12];
  assign CLBLM_R_X7Y120_SLICE_X9Y120_CQ = \ram.di [13];
  assign CLBLM_R_X7Y120_SLICE_X9Y120_DQ = \ram.di [14];
  assign CLBLM_R_X7Y120_SLICE_X9Y120_AMUX = \ram.di [9];
  assign CLBLM_R_X7Y120_SLICE_X9Y120_BMUX = \ram.di [10];
  assign CLBLM_R_X7Y120_SLICE_X9Y120_CMUX = \ram.di [15];
  assign CLBLM_R_X7Y120_SLICE_X9Y120_DMUX = \ram.di [8];
  assign CLBLM_R_X7Y121_SLICE_X8Y121_DQ = \wren ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_BO5 = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2663 ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_AO5 = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2661 ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_BO5 = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2667 ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_AO5 = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2657 ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C5Q = \wraddr [4];
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D5Q = \wraddr [1];
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A5Q = \ram.di [1];
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B5Q = \ram.di [2];
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C5Q = \ram.di [7];
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D5Q = \ram.di [0];
  assign CLBLM_R_X7Y119_SLICE_X9Y119_BO5 = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2665 ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_AO5 = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2659 ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_DO6 = \$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1517 ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_BO6 = \$abc$2590$auto$rtlil.cc:2282:AndGate$1870 ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_BO5 = \$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1522 ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_AO6 = \$techmap2616$abc$2590$lut$auto$opt_dff.cc:242:make_patterns_logic$1522.A [1];
  assign CLBLM_R_X7Y120_SLICE_X8Y120_AO5 = \$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1525 ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C5Q = \wraddr [9];
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D5Q = \wraddr [0];
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A5Q = \ram.di [9];
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B5Q = \ram.di [10];
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C5Q = \ram.di [15];
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D5Q = \ram.di [8];
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A = CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B = CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C = CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D = CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_CMUX = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_DMUX = CLBLM_L_X8Y120_SLICE_X10Y120_D5Q;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C = CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D = CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_CMUX = CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_DMUX = CLBLM_L_X8Y120_SLICE_X11Y120_D5Q;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A = CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B = CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C = CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_AMUX = CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_BMUX = CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_CMUX = CLBLM_R_X5Y119_SLICE_X6Y119_C5Q;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_DMUX = CLBLM_R_X5Y119_SLICE_X6Y119_D5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A = CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_AMUX = CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_BMUX = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_CMUX = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_DMUX = CLBLM_R_X5Y120_SLICE_X6Y120_D5Q;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A = CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B = CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A = CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B = CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C = CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D = CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_AMUX = CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_BMUX = CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_CMUX = CLBLM_R_X5Y121_SLICE_X6Y121_C5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_DMUX = CLBLM_R_X5Y121_SLICE_X6Y121_D5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A = CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C = CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_AMUX = CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_BMUX = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_CMUX = CLBLM_R_X5Y121_SLICE_X7Y121_C5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_DMUX = CLBLM_R_X5Y121_SLICE_X7Y121_D5Q;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_AMUX = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_BMUX = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_CMUX = CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_DMUX = CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A = CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B = CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D = CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_CMUX = CLBLM_R_X7Y119_SLICE_X9Y119_C5Q;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_DMUX = CLBLM_R_X7Y119_SLICE_X9Y119_D5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A = CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B = CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A = CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A = CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B = CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_OQ = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_TQ = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_OQ = CLBLM_R_X5Y119_SLICE_X6Y119_C5Q;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_TQ = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_OQ = CLBLM_R_X5Y121_SLICE_X7Y121_C5Q;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_TQ = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_OQ = CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_TQ = 1'b1;
  assign LIOI3_X0Y5_ILOGIC_X0Y6_O = LIOB33_X0Y5_IOB_X0Y6_I;
  assign LIOI3_X0Y5_ILOGIC_X0Y5_O = LIOB33_X0Y5_IOB_X0Y5_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_O = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y9_O = LIOB33_X0Y9_IOB_X0Y9_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_O = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_O = LIOB33_X0Y11_IOB_X0Y11_I;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_OQ = CLBLM_R_X5Y121_SLICE_X7Y121_D5Q;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_TQ = 1'b1;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_OQ = CLBLM_R_X5Y121_SLICE_X6Y121_C5Q;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_O = LIOB33_X0Y7_IOB_X0Y8_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_O = LIOB33_X0Y7_IOB_X0Y7_I;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_OQ = CLBLM_R_X5Y119_SLICE_X6Y119_D5Q;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_OQ = CLBLM_R_X5Y121_SLICE_X6Y121_D5Q;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ = CLBLM_R_X5Y120_SLICE_X6Y120_D5Q;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_TQ = 1'b1;
  assign RIOI3_X43Y25_ILOGIC_X1Y26_O = RIOB33_X43Y25_IOB_X1Y26_I;
  assign RIOI3_X43Y39_ILOGIC_X1Y40_O = RIOB33_X43Y39_IOB_X1Y40_I;
  assign RIOI3_X43Y39_ILOGIC_X1Y39_O = RIOB33_X43Y39_IOB_X1Y39_I;
  assign RIOI3_X43Y45_ILOGIC_X1Y46_O = RIOB33_X43Y45_IOB_X1Y46_I;
  assign RIOI3_X43Y45_ILOGIC_X1Y45_O = RIOB33_X43Y45_IOB_X1Y45_I;
  assign RIOI3_X43Y47_ILOGIC_X1Y48_O = RIOB33_X43Y47_IOB_X1Y48_I;
  assign RIOI3_X43Y47_ILOGIC_X1Y47_O = RIOB33_X43Y47_IOB_X1Y47_I;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_OQ = CLBLM_R_X7Y119_SLICE_X9Y119_C5Q;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_TQ = 1'b1;
  assign RIOI3_X43Y75_OLOGIC_X1Y76_OQ = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign RIOI3_X43Y75_OLOGIC_X1Y76_TQ = 1'b1;
  assign RIOI3_X43Y75_OLOGIC_X1Y75_OQ = CLBLM_L_X8Y120_SLICE_X10Y120_D5Q;
  assign RIOI3_X43Y75_OLOGIC_X1Y75_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_OQ = CLBLM_R_X7Y119_SLICE_X9Y119_D5Q;
  assign RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y44_O = RIOB33_X43Y43_IOB_X1Y44_I;
  assign RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y43_O = RIOB33_X43Y43_IOB_X1Y43_I;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_OQ = CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_OQ = CLBLM_L_X8Y120_SLICE_X11Y120_D5Q;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_OQ = CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  assign RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_TQ = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D2 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D3 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D4 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D5 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D6 = 1'b1;
  assign CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_CE = 1'b1;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_D1 = CLBLM_R_X5Y119_SLICE_X6Y119_D5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_DX = CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_T1 = 1'b1;
  assign LIOB33_X0Y1_IOB_X0Y2_O = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign LIOB33_X0Y1_IOB_X0Y1_O = CLBLM_R_X5Y119_SLICE_X6Y119_C5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A1 = \wraddr [3];
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A2 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A3 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A4 = \ram.di [3];
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A5 = CLBLM_R_X5Y121_SLICE_X6Y121_D5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A6 = \ram.do [3];
  assign LIOI3_X0Y9_ILOGIC_X0Y10_D = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y9_D = LIOB33_X0Y9_IOB_X0Y9_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B2 = \wraddr [6];
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B3 = \ram.di [6];
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B4 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B5 = CLBLM_R_X5Y121_SLICE_X6Y121_C5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B6 = \ram.do [6];
  assign RIOI3_X43Y45_ILOGIC_X1Y46_D = RIOB33_X43Y45_IOB_X1Y46_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C2 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C3 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C4 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C5 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_T1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign RIOI3_X43Y45_ILOGIC_X1Y45_D = RIOB33_X43Y45_IOB_X1Y45_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_CX = CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D2 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D3 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D4 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D5 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_DX = CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR9 = \wraddr [5];
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_D1 = CLBLM_L_X8Y120_SLICE_X11Y120_D5Q;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR12 = \wraddr [8];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR13 = \wraddr [9];
  assign RIOI3_X43Y47_ILOGIC_X1Y48_D = RIOB33_X43Y47_IOB_X1Y48_I;
  assign RIOI3_X43Y47_ILOGIC_X1Y47_D = RIOB33_X43Y47_IOB_X1Y47_I;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBTIEHIGH0 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A1 = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBTIEHIGH1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B1 = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR1 = 1'b0;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_DX = CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A6 = 1'b1;
  assign RIOI3_X43Y75_OLOGIC_X1Y76_D1 = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B6 = 1'b1;
  assign RIOI3_X43Y75_OLOGIC_X1Y76_T1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_CE = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOB33_SING_X0Y0_IOB_X0Y0_O = CLBLM_R_X5Y121_SLICE_X6Y121_C5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign RIOI3_X43Y75_OLOGIC_X1Y75_D1 = CLBLM_L_X8Y120_SLICE_X10Y120_D5Q;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_D1 = CLBLM_R_X5Y121_SLICE_X6Y121_C5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D6 = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_WRCLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign RIOI3_X43Y75_OLOGIC_X1Y75_T1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_DX = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_SR = \$abc$2590$auto$rtlil.cc:2282:AndGate$1870 ;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIADI0 = 1'b0;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y44_D = RIOB33_X43Y43_IOB_X1Y44_I;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIADI1 = 1'b0;
  assign RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y43_D = RIOB33_X43Y43_IOB_X1Y43_I;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIADI2 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIADI3 = 1'b0;
  assign LIOB33_X0Y17_IOB_X0Y18_O = CLBLM_R_X5Y121_SLICE_X7Y121_D5Q;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIADI7 = 1'b0;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_AX = LIOB33_X0Y9_IOB_X0Y9_I;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIADI12 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIADI13 = 1'b0;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_D1 = CLBLM_R_X5Y119_SLICE_X6Y119_C5Q;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIADI14 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIADI15 = 1'b0;
  assign RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_D1 = CLBLM_R_X7Y119_SLICE_X9Y119_D5Q;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI0 = \ram.di [0];
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B4 = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI1 = \ram.di [1];
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B5 = LIOB33_X0Y9_IOB_X0Y10_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign LIOB33_X0Y3_IOB_X0Y3_O = CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  assign LIOB33_X0Y3_IOB_X0Y4_O = CLBLM_R_X5Y121_SLICE_X7Y121_C5Q;
  assign LIOI3_X0Y5_ILOGIC_X0Y6_D = LIOB33_X0Y5_IOB_X0Y6_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B6 = 1'b1;
  assign LIOI3_X0Y5_ILOGIC_X0Y5_D = LIOB33_X0Y5_IOB_X0Y5_I;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_T1 = 1'b1;
  assign RIOB33_X43Y87_IOB_X1Y87_O = CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_D1 = CLBLM_R_X5Y121_SLICE_X6Y121_D5Q;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_BX = LIOB33_X0Y7_IOB_X0Y7_I;
  assign RIOB33_X43Y61_IOB_X1Y61_O = CLBLM_R_X7Y119_SLICE_X9Y119_C5Q;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_T1 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_T1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_CE = \$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1522 ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B6 = 1'b1;
  assign CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_I = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_D1 = CLBLM_R_X5Y121_SLICE_X7Y121_C5Q;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_D1 = CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C5 = LIOB33_X0Y9_IOB_X0Y10_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_CE = \$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1525 ;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR0 = 1'b0;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR1 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR2 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR3 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR4 = \wraddr [0];
  assign CLBLM_R_X5Y119_SLICE_X7Y119_CX = LIOB33_X0Y7_IOB_X0Y7_I;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR5 = \wraddr [1];
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D2 = LIOB33_X0Y9_IOB_X0Y9_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D6 = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR6 = \wraddr [2];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR7 = \wraddr [3];
  assign CLBLM_R_X5Y119_SLICE_X7Y119_DX = LIOB33_X0Y11_IOB_X0Y12_I;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR8 = \wraddr [4];
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D1 = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR10 = \wraddr [6];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRARDADDR11 = \wraddr [7];
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A1 = \ram.di [2];
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A2 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRATIEHIGH0 = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRATIEHIGH1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A5 = CLBLM_R_X5Y119_SLICE_X6Y119_D5Q;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A6 = \ram.do [2];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR0 = 1'b0;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D3 = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR2 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR3 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR4 = \wraddr [0];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR5 = \wraddr [1];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR6 = \wraddr [2];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR7 = \wraddr [3];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR8 = \wraddr [4];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR9 = \wraddr [5];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR10 = \wraddr [6];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR11 = \wraddr [7];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR12 = \wraddr [8];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_ADDRBWRADDR13 = \wraddr [9];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_RDCLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C6 = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIADI4 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIADI5 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIADI6 = 1'b0;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIADI8 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIADI9 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIADI10 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIADI11 = 1'b0;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_CX = CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_DX = LIOB33_X0Y11_IOB_X0Y11_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D4 = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI2 = \ram.di [2];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI3 = \ram.di [3];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI4 = \ram.di [4];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI5 = \ram.di [5];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI6 = \ram.di [6];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI7 = \ram.di [7];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI8 = \ram.di [9];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI9 = \ram.di [10];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI10 = \ram.di [11];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI11 = \ram.di [12];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI12 = \ram.di [13];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI13 = \ram.di [14];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI14 = \ram.di [15];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIBDI15 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIPADIP0 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIPADIP1 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIPBDIP0 = \ram.di [8];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_DIPBDIP1 = 1'b0;
  assign LIOB33_X0Y19_IOB_X0Y20_O = CLBLM_R_X5Y119_SLICE_X6Y119_D5Q;
  assign LIOB33_X0Y19_IOB_X0Y19_O = CLBLM_R_X5Y121_SLICE_X6Y121_D5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A6 = \ram.do [1];
  assign BRAM_L_X6Y120_RAMB18_X0Y48_RDEN = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_WREN = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A1 = \ram.di [11];
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A2 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A3 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A4 = \ram.do [11];
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A5 = CLBLM_R_X7Y119_SLICE_X9Y119_D5Q;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A6 = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_REGCE = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_REGCEB = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_RDRCLK = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_REGCLKB = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_RST = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_RSTRAMB = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_RSTREG = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_RSTREGB = 1'b1;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_WEA0 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_WEA1 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_WEA2 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_WEA3 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_WEBWE0 = \wren ;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_WEBWE1 = \wren ;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_WEBWE2 = \wren ;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_WEBWE3 = \wren ;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_WEBWE4 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_WEBWE5 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_WEBWE6 = 1'b0;
  assign BRAM_L_X6Y120_RAMB18_X0Y48_WEBWE7 = 1'b0;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B2 = \wraddr [8];
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B4 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_CX = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2665 ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_DX = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2659 ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A1 = \wraddr [0];
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A2 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A3 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A4 = \ram.di [0];
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A5 = CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A6 = \ram.do [0];
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B2 = \ram.di [9];
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B3 = \wraddr [9];
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B4 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B5 = CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B6 = \ram.do [9];
  assign RIOI3_X43Y61_OLOGIC_X1Y61_D1 = CLBLM_R_X7Y119_SLICE_X9Y119_C5Q;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C6 = 1'b1;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_T1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_CX = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_DX = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_T1 = 1'b1;
  assign RIOB33_X43Y75_IOB_X1Y76_O = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign RIOB33_X43Y75_IOB_X1Y75_O = CLBLM_L_X8Y120_SLICE_X10Y120_D5Q;
  assign RIOB33_X43Y37_IOB_X1Y38_O = CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  assign RIOB33_X43Y37_IOB_X1Y37_O = CLBLM_L_X8Y120_SLICE_X11Y120_D5Q;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_D1 = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D2 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_T1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A2 = LIOB33_X0Y11_IOB_X0Y12_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A1 = \ram.di [10];
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A2 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A3 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A4 = \ram.do [10];
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A5 = CLBLM_L_X8Y120_SLICE_X11Y120_D5Q;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B1 = \ram.do [15];
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B2 = CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B3 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B4 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B5 = \ram.di [15];
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B2 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C1 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C2 = LIOB33_X0Y7_IOB_X0Y8_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_CX = LIOB33_X0Y5_IOB_X0Y6_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_CX = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2667 ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D2 = LIOB33_X0Y5_IOB_X0Y5_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_DX = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2657 ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A1 = \ram.di [1];
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A2 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A1 = \ram.di [12];
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A2 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A3 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A4 = \ram.do [12];
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A5 = CLBLM_L_X8Y120_SLICE_X10Y120_D5Q;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A3 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A4 = \wraddr [1];
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A5 = CLBLM_R_X5Y120_SLICE_X6Y120_D5Q;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B1 = \ram.do [13];
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B2 = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B5 = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B6 = \ram.do [8];
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B3 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B4 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B5 = \ram.di [13];
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B3 = \ram.di [8];
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C1 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_CX = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2663 ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_CX = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D1 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_DX = CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_DX = \$abc$4086$auto$xilinx_dffopt.cc:347:execute$2661 ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_D = LIOB33_X0Y7_IOB_X0Y8_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_D = LIOB33_X0Y7_IOB_X0Y7_I;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D1 = CLBLM_R_X5Y120_SLICE_X6Y120_D5Q;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_D = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_T1 = 1'b1;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_D = LIOB33_X0Y11_IOB_X0Y11_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A2 = LIOB33_X0Y11_IOB_X0Y12_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A6 = 1'b1;
  assign RIOB33_X43Y31_IOB_X1Y32_O = CLBLM_R_X7Y119_SLICE_X9Y119_D5Q;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_AX = LIOB33_X0Y9_IOB_X0Y9_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B5 = LIOB33_X0Y9_IOB_X0Y10_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_BX = LIOB33_X0Y7_IOB_X0Y7_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C2 = LIOB33_X0Y7_IOB_X0Y8_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_CE = \$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1517 ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_CX = LIOB33_X0Y5_IOB_X0Y6_I;
  assign RIOI3_X43Y25_ILOGIC_X1Y26_D = RIOB33_X43Y25_IOB_X1Y26_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D2 = LIOB33_X0Y5_IOB_X0Y5_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D6 = 1'b1;
  assign LIOB33_X0Y43_IOB_X0Y43_O = CLBLM_R_X5Y120_SLICE_X6Y120_D5Q;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_DX = LIOB33_X0Y11_IOB_X0Y11_I;
  assign RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_D1 = CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A1 = RIOB33_X43Y39_IOB_X1Y39_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A2 = \$techmap2616$abc$2590$lut$auto$opt_dff.cc:242:make_patterns_logic$1522.A [1];
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A4 = RIOB33_X43Y45_IOB_X1Y46_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A5 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A6 = 1'b1;
  assign RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_T1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_AX = LIOB33_X0Y7_IOB_X0Y8_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B1 = RIOB33_X43Y45_IOB_X1Y46_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B2 = RIOB33_X43Y39_IOB_X1Y39_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B3 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B5 = \$techmap2616$abc$2590$lut$auto$opt_dff.cc:242:make_patterns_logic$1522.A [1];
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B6 = 1'b1;
  assign LIOB33_X0Y111_IOB_X0Y111_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_T1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_BX = LIOB33_X0Y5_IOB_X0Y5_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C4 = LIOB33_X0Y5_IOB_X0Y6_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_CE = \$abc$2590$auto$opt_dff.cc:242:make_patterns_logic$1525 ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B1 = \ram.do [14];
  assign CLBLM_R_X7Y120_SLICE_X8Y120_CX = RIOB33_X43Y45_IOB_X1Y45_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B2 = CLBLM_R_X7Y119_SLICE_X9Y119_C5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D1 = RIOB33_X43Y45_IOB_X1Y46_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D2 = RIOB33_X43Y39_IOB_X1Y39_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D3 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B3 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D5 = RIOB33_X43Y39_IOB_X1Y40_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B4 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_DX = LIOB33_X0Y11_IOB_X0Y11_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B5 = \ram.di [14];
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B6 = 1'b1;
  assign RIOI3_X43Y39_ILOGIC_X1Y40_D = RIOB33_X43Y39_IOB_X1Y40_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A3 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign RIOI3_X43Y39_ILOGIC_X1Y39_D = RIOB33_X43Y39_IOB_X1Y39_I;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_D1 = CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A4 = \wraddr [2];
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I0 = RIOB33_X43Y25_IOB_X1Y26_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A1 = \ram.di [4];
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A2 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A3 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A4 = \wraddr [4];
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B2 = \wraddr [7];
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A5 = CLBLM_R_X5Y121_SLICE_X7Y121_D5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A6 = \ram.do [4];
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B3 = \ram.di [7];
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B2 = \wraddr [5];
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B3 = \ram.di [5];
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B4 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B4 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B5 = CLBLM_R_X5Y121_SLICE_X7Y121_C5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B6 = \ram.do [5];
  assign LIOI3_X0Y3_OLOGIC_X0Y3_T1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B5 = CLBLM_R_X5Y119_SLICE_X6Y119_C5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C2 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C3 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B6 = \ram.do [7];
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C5 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_CLK = CLK_HROW_TOP_R_X60Y130_BUFHCE_X0Y24_O;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_T1 = 1'b1;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_D1 = CLBLM_R_X5Y121_SLICE_X7Y121_D5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_CX = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
endmodule
